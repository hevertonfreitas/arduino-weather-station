PK   ��GW���Ք'  C�    cirkitFile.json�ے�8r�_eC�-v A���۱=s��	�c}�ݡ�Dj[�R[���;�ݍ��$��@���8l��_��_����~�������a��_ܒ�Y|j��/�ۿ�������[�c�|�������~��e�}״�]�f�Z�5��ˬw]��e����U۔�:/}Gf�gq�����
$Vb��Yڠ�z���/�>�7ۻ�뗟ww�~{�-\���ݎ�N~r;��O�w���aY:ڬ��f�um��~����de�Y_�TU�XVB�\���!U0K/�����?�&���)�&�*�e)f�*���R��Y�b�BАG~�D�~y�'i�%�D��M�Ky�Ki�#�D�M�D��M�D�N�D��N�D���c�X"P�c�X"P�{�خ�<۩�sW�]N�f+KU���˚ژ�7�h��7��C�]x�n���8d��ʛ+o��B��%��9K
ys ���@,�mys ���@,(�]i�D��w���BޕK
y�K
y�K
y�K
y�K
y�K����N�D���N�D���N�D���N�D� �c���N�D���N�D���N�D���N�D���N��Yzy�K
y�K
y�K
y�K
y�K
y�K
y�K
y�K
y�K
y�K�e!��b�@!��b�@!�����AGs:,�����GCadáU�m
�|�����Jj����<�����oTf7(�tW;���N��53�`0���LNNg�9��s��t��I"�vk;(a�N&�!l�C�5e�����&3U��|��Z(a�̲�ڮ��JGX:�����������,k��j��t���y��>}��{�P>��^���I:+����c����	���|<kl?p���#0�����`���3������	�G`>�c�8�����W���:�|��u`��3,��xE�~���G`>^K����X>��*�������|����������p�b���/X>�.U��/JD��~+���ܞ�\��ǂ�,��xI�~���G`>^�8���������~�|���`���,��x�$x�	8�����}���~�|���`���,��x�-�~�b�)b��%����jo
O4�ޔ�'Y��5Td�ݴYS��m��Za束�|f��0뉭�Ӄ<5p֓��,��x18�~��G`>^��8���������z�|���`���,�����~��`������g=X>�q�	���Y���|\"l?pփ�#0� ��6�8�8p��ά��Y�P����h�ք��R��M%˒OQ ^�z�|\�����G`>.��8����������z�|��rEX��3uf�b�4��ȭ	MN�<8a�����K��N��|��X`��&,�����~��	�G`>�E������|\El?p��#0����`��Ǖ����.X>�q�=�������|\-k����G`>�s�5��j�,ۃs,Ww�n�\�,�����F#��VofջayЙ��zμ|X�s���*ĳ�I���]{PF2x$�2�3/������l)S.��a�޹���U�Kd��\�lH'�\����?-zh�6�s�V�{����6=�{������kI�(zt��W������6\��ys�z}�����Q�ʈ�])�m�v%�m+�mћJ�W5��m����[]֛�׷��̹u��r�f�MY�f�Yc��R�.���˞t���^��u�\�n�uh+�U�.2jlcm���m��{�����t���'���F.��e����"4�To+��&�i'����8iK�����(RWNb��v���GX��2O�%?-�>x8{A��%V�S������>�.�N>�.��=�.�N�S����@��.E�=��va%�-z��'�+?���F���_{��a�\��v���IX���L���=s��2�fb�@B��J��{9�E�S�2�E�PO$�[!��?�dDET�l2ܬc�@B�{
"�����$d��(D�6.l��6��-��L�/1�b7��7J���&,~,���L�Y����(%��1�⸅�q���?x��p�o\�m}7��+d��q�P]^���QJ��(	b��q��(%��1�⸅�q���?zb�PJ���
b����G)q�>,���8J�����`q<��q��1��x��(%.�c��q��(%.�c��q��(%.:c���aq���8J�g9��`q���8J�K���`q���8J�gl��PJ\c����QJ\����QJ�f����QJ������QJ����,���xj�	�X�R�?mi��{l�^��/h�/τ��
�Y�gc��p�6B�TX�%� ��^c�u� c���
c5�a)*�*Ю����.�Ua,��J*���b�a+L���J#�KZ�U����J*�f9,uW�U��TX�rX�
��+����4\hWVRa�9�:�A�� l�BK:�<�YǶJY�RڥA�s�ul��y�В-�5ױ�N��BK:�<g^Ƕ:�
-�����jd6�CK:���AǶ:��
-���Z��dc*��C�kJtl����В-��ѱ�NV�BK:���GŶV'/S�%Z^��c[��L��thy͕�1�/bJ��t�2���Y��L��thy��m�L�G���h!F��ˬN^�BK:��&QǶ:y�
-����J���e*��C�kDul����В-�uձ�N^�BK:��fWgb�N^�BK:���XǶ:y�
-���j���e*��C�k�ul�4[Qi��N^6��O���e#����e�N^���e*��C�5tl����В-�Jб�N^�BK:�\�AǶ:y�
-��r�
���e*��C�58Tl�t�2Zҡ�Z":����ThI��k���V'/S�%Z��c[��L��th�F��m�V�)-%��˜N^6ܟ����-�q��Op:y�-Zi[�����e*��C�5�tl����В-עұ�N^�BK:����!F�T�P��1Z�t�2����В-�8ӱ�N^�BK:�\�MǶ:y�
-��r�9���e*��C˵�tl��L��th���mu�2Zҡ�Z�:����ThI��k2��V'/S�%Z�-�c[��L��th�F��m��e*��Coc,t�Z�,Ҷ:y�p�d�x�
-��Ʋ3�Ξ�t;Se�6��m�!*u�g����w��Ħ�3U&�[�T��G=S�XA:�Jz��D��^r^��7}�;c�N"s��έ��L���+3Q�}�ƅ���+3Q}�̓�M^K�^�ŵ7&o$2��	�S�TΕ�x��^�se���lW^"�{qM�Y�$2O^L�I�㾆�M����5��\��^\��&�L�+ʜ[��*7m�ڔm֛�1�r�&I�r�JR��>�k�'���f����Ye�"��6ֶ����]�T.�%I�]��ԛ�ܰØ�BEV�M�5ea]Qۦ�����%�Х~Z�
�.��I*�Rg�+�.'c���*s~�eMmL�[4��_�G략K�
]|F)*���;(�T�/��I*;'�T��$��]�$��=�$���$���A�יK�u�]j��d��:M&��Z��\Lo�d��_{��a�|84�nq��Uw�&5����þ�{8�����$d��!	�>�B�@B���"���>�$d�B2}k!	��e���L�JB�@B���bB$.j��6,n,p��̱c�a��n�o��9vy0L��M� �R2ǡZ,�,����q����QJ�8��a���qpX��8�R2�Q|,�[XG)���,�[XG)��,�[XG)��7L:��9,������	7��J����QJ\u
���9,������	�sXG)qU,�;XG)q,�;XG)q�nL7(���QJ\�����QJ\M ����QJ�z���=,���x�4�	�=,���xu.�	�u�y�=,���x%�	�=,���x��	�XG)�*1,��8>�4�W���z\�P%VRae]�F�	!�`%V��V�U�v�`%V�����U�v�`%֐w��5*���+���~��]��.h��
k裨�5*���+���eT��
��+���eT��
��+���eT��
��+���`��@'�R�%Z�۬c[��K)��ɻH'�"��K��thy���mu�/Zҡ�9�:����ThI������V'S�%Z^àc[�LL��thy-��mu�1Zҡ�5%:����ThI������V'+S�%Z^��aA'/S�%Z^��c[��L��thy͕�m���)}��ˬN^fu�2Zҡ�5p:����ThI������V'/S�%Z^��c[��L��thym��mu�2Zҡ�5�:����ThI��׺��V'/S�%Z^��31I'/S�%Z^{�c[��L��thy��mu�2Zҡ��:�U���4]Q'/�u�\'/S�%Z^��c[��L��th�ƀ�mu�2Zҡ�Z	:����ThI��k>��V'/S�%Z�]�c[��L��th���m�N^�BK:�\KDǶ:y�
-��rM���e*��C˵]tl����В-רѱ��J2��d:y���˜N^�BK:�\3HǶ:y�
-��r�#���e*��C�5�tl����В-עұ�N^�BK:�\SKŶ^'/S�%Z��c[��L��th�ƙ�mu�2Zҡ�Zm:����ThI��k���V'/S�%Z���c[�*Je>t�2���y��L��th����mu�2Zҡ嚌:����ThI��kK��V'/S�%Z���b�B'/S�%Z���c[��L��th�f��mu�2ZJ�}�+�t�Y����̭�&[9��ʶ��j��B�c���L��ڴ3U&���T���=Se���L��Z�3U&�[�T��G=Se���L����s�����u����V�+���L��`|xj�й2/�ڌs�(c�xj�ʹ2/��r�Ƌ�v\�+���}綺/��=�U�.�M���W�9�γUn�l�)ڬ7+c��^M�
�����r�}*L�:O.[��:sM���EF�m�m��e�$�\�K��E�t��7e�a�1A�����6k�º��MUW��(I��%�`���NR�8���r26[Y�2�W]���d��EӬ��u�`����MQ�l����MQ�X�b���r�QJR��&%�\l��T.�Hi^r^��^��d0�{9;H�y��_o¿�zX�ww��r����%s��e�����u�.���ݾ��������he0����z#��oHBgHDjl�7dWl�-����`��U��O�
SZ�`�j�G��5��~b&�d>ڹ[�Pd�G(|�PQ��\�x��	�pٷ��P�4���hlU�ӹl<v��2(�.����r�(A�b���3�C-�ia�7�Q,A�+X#�Da�~���;��E�V�d%�]�~�$�]�~�H~�X|����v?�$��o�����2�����a�z98���84�GsP��o>ta�`��| �l� �*�0��4GCЀ�A�a���F�(4���x��N�&d���J:q�Ɉ��=�$'��/�	��L�	��h��=�$'�=�!�CPr�H��H: pV�� 	=<@��R��U � A<tŃW!�=n�wˇCs��/���l����n��m�_$q�g�,%������&�K�~*�9�G�*Q�(��c('���PN������70M.��r�Bn����
)���w(�K�~ޢ�B,a���1j�lI	�a�S7���J��*�0�ɣR@%@ �k���6) � ��5�qy��O- ��5�q����y�z! �ڸ�J���D�~��Z�|- ��5�qI��|- ��5�qQ��|- ��5�qY��C�a��R����:�rޤ��9�3+��ͯ �x��\�7Up �i��rެ���O��	�O ��5xs b�1�
��O������O��q �O ��5�3��C�����x��T��E��x��T��Ŧ�x��T��E��x��T���q�xZ �\��� 8 � ��XC<E:�N<�
��K�|4YKM��қ�lp�*�����H�Qs
��F�y�I��F�8= �YFۤ�� ����/d2`�E{���G`����E���C.�},.Ÿ�ۏv8��A��G`>��v1��A��#0�YF;��� �����,��Hpz�a��ǳ'ѽ�(;�v����&䙟h�Sx΂%�Y�h�0!�	y�-چ��LHhB�-��!:A��g:�m�����Є<KmCtf&$4!�0G����		Mȳ��6Dg(`BB��~��Y
��Є�*lC��S���&�h��0!�	�X痆��1&�PA�-��Xt�&$4�iU4����ܢ�+,��bb`��Y�Eg1`BB�r'��Y��Є�TmCt&$4!/3C��ŀ		M�K��6Dg1`BB��>��t&$4!/MD��ŀ		M��*�6D�-`BB�P��S��s��i˰,j�e�8��,�����R����ŀ		Mȋ��6Dg1`BB�i��Y��Є��mCt&$4!/LG��ŀ		Mȋ��6t�,LHhB.��!:�����m��b���&�Bh��0!�	��چ�E-�U-�<š���Q�<�5``�Z J
-�9��x):�rY����0!�	��
چ�,LHhB.��!:���tG�J���I8eL#�R���Nj���&�Bh��0!�	�چ�LHhB�䄶!:����P�m���&$4!W�B����		M�տ�6D�-`BBr�2��i��Є\umCt�&$4!W�۰@|�0�$2�Ԅ�N
t�1&E�-ýE�g$�������UF5�n�+�>��8�������G�����9���d?Ө"���J�3���ۑl2��lbo��+ś4�v��7��I&�@n�@T�x���g���
Du{�o=�&ڑ^)�]iԍw�+ ��x����4�m�]�z�ݴ#=��رS[I�w�+pƋ���]h}E�s�<[��V����z�
��.I�K��K�t��w�0]�<�l�6��5��*S5������6��?��3��t����So�r�`��Td�ݴYS��m��Z�Q�t�L9��*������$���:��H��~�E�VIr��i"�&ɍt�&��Ir#�b�9O�y�@.N�:Irg�_Iן�}%]��t��!�cמj���bߞj���b�j���b�j���F�{*,'��w��z�x�ٶ��n~�aq�e��yXܾ_�M���a����5���q�g�>N���q}`��I�W������V{���ҽ�X������|��+,_���C�1�dB��S����E)mǸ���燲�������;�s^� a��^?�#Y�'��Z��FE��� b8'�;�u]����?�jom��7�	)��w�::1ayB(z;�Po�8���Sh�K�;�	�w�K��&^��LJ7\[��:�Hå�M5A�y�hp9��j'�P��tLc�hҒN���K^O��N���E1�T����U;�0�H�Z�M!�����1])�~<�i&�{bF�b�M���:�"³�>1���8�>q8A�!��x��ːT�8��.���7Y�����kV�'�f���v�o��O�s�#�t��C�鐋��C>>T<*�C�ӡ2>d���P�t(�UO���P�t��ѳ5(6��#�=3RIϐSҳ)6$=�bKҳ%)6%=��b[ҳU(6=��b��g���.��.6��}yv�]�]¿_m�B�|�l�7�������PR�,������[���~�Oڍ|y�m���.?��>�Ks౯/��~��>w�ö��|���_�`���~{���}��7�Y���=���MV��~���E���O�_�z��Awq�i��p���}��]�u/�w����w������j�7������ ޞ��d�>n�w ��Z��a�vx�����toLzc�}���LL˴?���ەw&�J�MV:��cWY�
˗�t��n{�ph���k�Fho��6<��H�x������w���|�YS�{�Z�7y�?ބۨ���r�,���׸�k��kh�3uM9u�Oi��+�����燗<<f�bL[��%7�yw�\�+NO���rJ;����?�P�yTCc��WR�y>Q�%��D��Fϫ"�=-v���b=-v��g��M�΋]7>�c>�k{�������������;Z?i�W���m6����O?ܷ�|M��o%���KOv�7�>Z�ro��M���f]f�w�̮V�������V�k���C����!>�o
oؓrw�$�r ���/GȎ�ʑ��{����#m�)���ׇ���GJ��|ǟ�f��Dǿ<����	��c>�H�<����x�d�Ma�w���������3m�|��ˬެ����*߄���\���#M�6��H��Y�7�KC�#_?�<	�(_"�)�+���k����L흫^�j[�se� ���\H)��3���|cBSX�Y�o��hu����&��wSW��zM9��w7<��eU��q�:��c��'?��2��ᒯ.���j[eɆ.؏r�&2���]]�mz
����*��]:eiJ�d��&��;�;���'��UW�����]��W�f��Fg�f��2���S'L�Ο������\(���T�w�| s�+_��k���I��Iμ����/��������x/���_��dgz�|���s"�{�o{�>�,�S��ק�������~ٶ�O,@�zgÛ���m����7�.����:�����<��Y���^2������߷�/�ܭof�|/��n�aq�a�O�ϗ~X�|o@�?������]=����)���^z���7$j��W=�ϻ����������Ç��u�#�[u�������y�ks������g܌��u����?�������f{�t��7���k�94������4�sQU��;�9�L�3��!ǣ�g�vv��mR�9=�U����ƽ"d'�(�z����8��l��.{x\e��ɔKs�+�B�B�il�������?�44���&~r�PIg�N|uKw��B`@�f�9b������뚾L�L�	��5�f�&�ܬ&I� N�F��:�Mr��Y>-$8�t2�V_7� �:}�k�a�׍��S'��9m�WS]8��l^����j\B qJk[��}�������=~��#�?�uz�ᚖ����>�ׯ�����pg>���$��o$'�{xV�s�7~x��H;��m`��W�6Ѩ���]g����Ps�Y��3X�����i� ��4zp��(Fuy�ic�CKl�Θ�C��ѹ��܅:���'��q�x�G���NG|�ч>��);���x��'���:1�عuCPKFL[}�v��b�5.��`)�s��%�4�N�W��8�U^U~p��܈ē^&O<�������y��U��ww�+�_�j3�7����1;�H;K����.�:ŵ}�tV����u���/��뜞UU�;�'�zq���&zjCgM�m6]�D�\%��I�_��f|���:���A���ʍ�]~�Y�O�����5��U���㪡�qU��_���y���଩��i7(�|܁���R��Y�~���>�\Ŋ<��y��y��;=k�-+lJ�W\5�����칎��J � e�m��.@���NϚ
=�O=�,;�:�bI'}� E�O=�"�>9xj�8�L?��£�9k"S�.%�����9l�6(��vx�6�;�y(�}�5�ryJi�gMdtCwM��꼄��[`7���t���u��G5����GOr����8�:#�V@ϸ��_�Dv?��'��W�>'�/jj�z�������t�_���qzR6>4t\�6󬉖�������Oٮ<��
����X?3W�Y�NO��?���,�5��~r{w���_�C��6w�=Zp���?��ӵi����v?�p�~z����u��PK   ��GW���Ք'  C�            ��    cirkitFile.jsonPK      =   �'    