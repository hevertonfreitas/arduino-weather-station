PK   W�dWi���/  ��    cirkitFile.json�[�丱��A��R���.�f�?��`��>�4�L�S؞�ުj�����T�-E�����`���)*�S0d������p�;����7w�W)\_������j�������v���x������__�j?���]�g��75G_���ʷ���C�V�c�tׄ��.�������/�@b	Q��A*��l��z������꾿�̾���s���x�Õ�u��u����~�rw;�>�O�nl�[��!���۱j����6ԻV����^lR	f�^-�v��P�A�:�X�R	f׈�L4n)�T��ub��(C���"���;�:\���B�~��"�����B���"�����B�nS,"
�;N��(D�:�"bgO�;�""��w�ED
q��u��a[�<M782��[j+�C�w�T��u��	]�����p�U�}W+o��9����@,"Rț��H!o�""��9�����9����@,"RȻ�b�Bޕ���XD���N��H!��b�B�;�""��w�ED
���0;/��b�B�;�""��w�ED
�����!`���r�))�S,"R�}�XD���N��H!��bf�S,"R�}�XD���N��H!��b�B�;�""��w�ED
����r�))�S,"R�}�X���r�))�S,"R�}g&b���9��`�\�,�����C������W�ʃ��T�Y��,�����;��LoP:��.6� T�-��%+�`0�J��&NNgvk��;(a�b��՝��JGX���s݅�+�da�LU�w���d������V�#,��5X�5X�A�Kgv-Vw-VwP:�ҙ]��]�����ti,�O�E/�^8���|i/X�A���c����	���|i�4X��G`����?p���#0_Z���?O`>�5�`��#,���� ���Q���|i_X���G`��#�?p��#0_�K�՟�X>�]0`���,����7����
zz=�_,8|����G`��J�e��s�¹�����	��~,8����/m)��`�̗6Á��~�|�K����G?X>��`���,����I�p��#0_��	�8����/mW��`�̗6ڂ��^!�^"_\ֿ��&�Do��iƴ��T���j�x������l�v��#o�N���QO��<H����z�|�K����G=X>�m�`���,���|���Q���|)u X��G`��� �?�z�|�K���G=X>�D`���,��R����Q���|)�X�1��1��Ã�������eQ(�_�^M��,4�XU�(�b��˗Ѐ��`�̗R���z�|�KI��G=X>�tEX��w�lt��e�W��W�
0p���#0_�.�8`���/���0a�̗2z����|�K����O�`�̗����]�|�K�����.X>��u`��C,��R�=�������|)[ V5x��G`���7j&���Y �g������؛�[��6U׌�2��w�SwI�n�j)1$�쳰�r3�fa¾1ߍe�c�s�͓�n�}�Mt���4�o��>ޜ�R-k�指2�ه, �'/�x�<���de�����Y��~
�OI�-�-9H�L/��t��ŏUZvx����9÷�/�`����?ϰ���NҬ��n:���GѣI���޺���mE�����|[�~k�ix�wE����˟M�g��g�lF�H��d��m��ܢvM7�!�-U�\�w�X�Ǧ��0��Y��^��n/��>�����6T���z�[{tc�wޝu{��Y��ߝ��E�~��D�B@�rמ�"Tj����!
�E�.�?�5Y���	P��4_�%@9��\tf���2K�$���<_�!@	-�Rg���r�ú��n/G<���a>�)�{-� ���ۅ�<��p���g��x+��I����%,�q�|D��E��4�a��&�6����?���wGk��0�cmcK��z�(v/}�'�B�Ҁ�ɥ������ɥ��ɥ����R�zr�g=�4����+5��G��x�.30�d�<����|.s�M���b�8���"[(}�Lg%xr�g:h��K_=�Q<���3b��K#�̦A��Ҹ"�i�8�Rׅ�6H]�0ۆO�N��=��w���>�"	ã"���Lޞ��<O� �?�$(����Or"�"r� 2�ndDE�Q��]������G/#
(��#� �ZH�I��$ȤV
Cd���"q^�a~�@��`��4�b��n�9o�$3�s��`��`%�L��@L0N0'��d�EN &��0?��d�eQ &\����q;y�q��B&����0?na~%�L��@L0?na~%�L��@L0?na~%�L��0L(IfZ�b��q돣$���0&�w��8JRJ8c��q��(I)1.�	��̏�$��0&��0?����`~���8JRJ�	c���a~���8JRZ�
c��q��(I)}�	��=̏�$��(&���������Q�R�.̏�GIJ��`L0?`~%)�=�1��x��q�������5̏�$���0&��a~�$i�2�yz���{��)c��h�8���TX�n�:S[�,@��%:�u��c��?�`�0V���I�K�U��TXcܥ��yU�4XI�5��T�:O��i�4Xi���y�U�T��j��
���Ӱ¥���J*�f7O�
�
ԫ+����<m+\*P�����y�Ё
-�Ц��:�U����.ڴF[G�:��
-�Ц��:�Չ�ThI�6���ѭN�BK:�i�n5"ҡ%ڴ�AG�:��
-�Ц�:�Չ�ThI�6�)�ѭND�BK:�io��nu�2ZҡM{|Ttku�2ZҡM{�tt���Вm�s�3!�4#�4%��Y�����e*��C�����6�t38*��DQ�N\fu�2ZҡM{ut���Вm�[��[��L��th�Q���e*��C�����V'.S�%ڴgWga�N\�BK:�iﱎnu�2ZҡM{�ut���Вm���[�ՊJ�u��y*����(��l��[�����eN'.S�%ڔc@G�:q�
-�Ц\	:�Չ�ThI�6�|�ѭN\�BK:�)w��nu�2ZҡM98Tt�u�2ZҡM�Dtt���Вmʉ��[��L��thSn���e*��C�r���Vi'��V2�����e��$A1�
--�B��G:����-Т�"u��y��L��thS'���e*��C�rQ��V'.S�%��Sk��u2z���-D	:qYЉ�ThI�6�8�ѭN\�BK:�)W��nu�2ZҡM9�tt���Вmʝ��[��2ZҡM9 ut���Вm�e��[��L��thSNF���e*��C�rK��V'.S�%ڔ#SE���|�
-�К�q�c���В�9;)i�y��OP�%��C��n7J)��z =DJ!��F)~���(�p��F)�����Qo�r� �%�QJ!��V�/�zO��v�1� s���z��)���*���}��	���*��}��'+��$^o��.�z��Ɋ�v���9Yq��C+��¥�%���X����q$b&+��h{��'+��%���\�q�\#q[����Y��]Ӎn�b�������������4ƽ1v�WÒ�aY�հ��~O��>����P��Uk���������~]/,)�zaIY��Лnl�1��R��Z;�����;۷]{z���i,)��OcI���j�ϒ��:#C�������ʇ�P��1U�m���`Bם���^8Rh��8R��O�OP�(ŭ��,)���7J	k?K�j׊%e�gŒ�ڱbIY�xVg�Zk�Zk�yb�Zk���Zk����'f5���3M��	�W�z_�G�W�`��h����V���@�TO��Q 婚���_����꾵������;������]�~YR����Q e�2a쏾��á�۱7�!��m��Ce�]ﬧ�8�z�Ē��*����K,)n-vcI�kVǒ־ ��z�kdIi�<KJ����tk����ڇ�Co��_'9�ǻ��c�8\}��U�����������p��` Af�R!D Af��!D Af� "� 3y#H��<�$�L^Bd&�!	2������%���S��q�8��s�0�M0Ǎ�dN!�	�	�Q��)��0��7�8J�9M�a�`>�`N%ɜ��0L0?na~%ɜ&1L��7�����Q��i������Q��if�����Q��i������Q��i6������q���GƄI�������q���������Q�R~9̏;�GIJ��`L0?�a~%)�ς1�����q����	Ƅ�������q���W�����Q�R̏{�GIJyC`S?0?`~%)婀1��x��q���Ƅ���Mo��x��q��������Q��~i̏�0?�����`~�����{m���h��-� ���J*�I��^�m�h��
��e{��R�z�`%V���j�����J*�1�R�k�R�VRa�� �f� �`%��GQ�k�J�VRa5�,�Z*P����jvY-�T�^5XI����Yh�@�j��
kZ��D\*��C��6��V)�R
�t�.�	�H'�R�%ڴ�\G�:ї
-�Ц5�:�Չ�ThI�6���ѭN�BK:�i��nu"1ZҡM{1tt���Вm�S��[��L��th����De*��C����L,��e*��C��*��V'.S�%ڴ�JG�J3bJSb:q�ՉˬN\�BK:�i��nu�2ZҡM{�tt���Вmړ��[��L��th��J���e*��C�����V'.S�%ڴ�UG�:q�
-�Ц=�:�t�2ZҡM{�ut���Вm�C��[��L��th�^p�*�VTZ���9�����e*��C�����V'.S�%ڔc@G�:q�
-�Ц\	:�Չ�ThI�6�|�ѭN\�BK:�)w��nu�2ZҡM98Tt�u�2ZҡM�Dtt���Вmʉ��[��L��thSn���e*��C�r���Vi'��V2�����e^'.S�%ڔ3HG�:q�
-�Ц�G:�Չ�ThI�6�p�ѭN\�BK:�)��nu�2ZҡM9�Ttt�2ZҡM��tt���Вm�q��[��L��thS�6���e*��C�r���V'.S�%ڔ;OG�JY>��|��eA'.:q�
-�Ц\�:�Չ�ThI�6�d�ѭN\�BK:�)���nu�2ZҡM92Ut[��e*��C�r}��V'.S�%ڔ�TG�:q�
-�h_ϊn<����Uo���0V{oǪ96�Gj���(d��(���v��B6ٍR
y�7J)d��(��+{��Bv�R
��7J)d��(���y�Ձ�c��C_����o�hխb0\:�t����	�*cť�8���`��N��*cť� ���Xq��ŭb0V\:�pk�����遯b����CK��W�9V���i<�{c�z��%ò�A���~O��>����P��Uk���������~]/,)�zaIY��Лnl�1��R��Z;�����;۷]��F,)�oĒ�y�՚fIYu�C�������ʇ�P��1U�m���`B�1�ˑ��]��u�r��k�#���V�%e�QbIYm�XRV�$����gu ��X�zt������'fՂk�L��jlB�U��W����0ؽ;Z�7�gIYo�8RV��%e���HY�$�L�z��U/s8�};��:��V��M�5c�̾���GZ���U{aIY���U{aIY���U{aIY������J,)����@���z���g���������ϫ��\_�|s?<�|��qws���?�W��^0(*����|���$�H�@�7$�wHDҒ�ߐm?&�Jaf�"� ��V�pw��Tie�T�|�R�w�g�ډ)��v��>l��B�!�PX�P��N�*|��q�<���P�i,�cA�Y-ɣ�l&��h�ؕ���$(B��o��Xa�@V'"s�D��y�� Ђ52K�����J�+�D,˴2�$+yv+{6I��Ȟm$ϮK�f�I�Y$O.T6shF��BU3�s$O.T4sH��F6�"yt-%�<���0��$O.t5��t�'3��k+%(��^�2W�"jZ�]昶h1ӧO�#���Ow������4��}��������͐�<r;�~hUQV��o>0a�O�+^>L�����6�
=��9ͱn4 |�{��a����7���I؄���(=�'
����d�@N��6�Ig��I��	��\��=� '�,�!�r�<��H:� 0V�� 	=� @��A �S � A:1�.�o1?!NS���r ᤅ@:w!'�Na�	�3r �ƻ �d^CN��ސIg9��Ɏ4�{�_on�v���p����w�x�{��}�9^}�E��N+�w��:�E�i���B,�L�7��Qs�"�r9��A99��חX��6��T�dPAU�U#a��2B
�3�R�E�i���B,��H}��"|-�ْ�7@�9m��r \*|�\�9m�r �(�\�9��r |)��\�9%:�r ���S�sJ�$�@t^z�A�p�6ￒ��j�v�%5�V-�8_p�r��J�p��|�2�)����|-���e�S�/!�\�9e�r ��tf�2�q� �{u�ά\F:����O�2��� �?u *���Mp ���S��t/��O=���e�c^��VĀ+��z�?��H+�  ��T.#�� �S�riᔜC.#�� �� �r�x6 ���?��H�~8 �4 ��\F:N
���O�2�1E �?��T.#-�p �i��lHS�T=;i&���϶a��UXz3�?$���$��lRޢ:���S�f�q۪ ��pq� |f�X������|1��/;�V��X>�mσ�/;qv��������
_?;k'b�X>�]v�,NDX>�]vf,NDX>�]v.,NDX>�Փ��vH��XBB���h�Cx̂%L�V�:D&`BB��h��0!�	�ja��
��Єi�3Z��^?�		M�Vi�u��L���&L+��:DG'`BB���h�#0!�	��~��Q
��ЄiWX���		M�vT�u��S���&��(��5D&�R��
:l��Ţ�0!�	��hbt��m�@�(&�j �Xt&$4a���!:��0m�B�ŀ		M����u��b���&L[��:DG1`BB��}��#�(LHh´5�Ct&$4a�V��!:l�0m	E�����igQF���ŴB����X�at��Q��Єi�1Z��(LHh´A�Ct&$4a�܍�!:��0mLG�ŀ		M�6Ճu��Q��Є)! Z��(LHh� �Ct&$4aJĀ�!:��0%�@������xt�2?(K�'<�L�RdA�L��=��1V��b��)-	�J�Q��Є)�
Z��(LHh�Ct&$4��`���+��I�dL�R����j���&L��:D5`BB�lHh��0!�	S&'��A��Є)Z���0!�	S-��a��Є)�Z��LHh��Ct�&$4aʺ��!:l�0e��FO��		M�+�Ej�e'5:lYv�,=`��1V���*���G�fU&9N3����v��Y�ō�g�f7޿pȌ�4��%�cg�Z7ޟ�Y�x��N�]��,��Vc[��\)?�It��t,�L��`���
�Ro ���$�����[ty����8��+�=�8kD|�Q;�g����U�Ԋ���
�3�Xљ�M.Ot
v�o���į�'Gm����ntCp-U�\�w�X�Ǧ��0�#�{����ӱa���7T�����p����P���+�mo�����{���?��w��M76͘�����Z;�����;۷]��}�����r�y�b�8���}���[�M782��[j+�C�w�T��u��	]��{*8+��\�T�,q]�Bk��P�Ɣ%n�*j��<�(uX��霱��oƺ�����w"�)�]j�y�r�.��<y�q��u��ܺK�:Oނy��2Kނ}�r�i��X�M������?���wGk���j�����P����%n�r��%n�n��%.�ZW0=���f]��X�:��c�[���p��v�Mu��|c��k�P�}�;�;��`w�Q9��� ��X���K\nw��%.������vW��X���X���X��0��Ͳ��Q`���;.|�<y�������U��q�x��x����'Լ���Uzɤ��ͦ-�_2�Tөz�kH�S�z�O�;u>�.��ћ�gS65�Sk;5�S�`�lL�=�dJ�L�gRΤ�X���#�b�o�Dh�7ƛ8�Ʋ��͌�������(�cw�p�V��d���c��]hf���'/DK��UѬ�LV��$yQQ*��\��K���p���x.8�^z�]��ZJ(��<�\N؜���� �ױk��js����O��2��-|�̱A�<�FN�I���dtTj��#���Ԝ��N0�UES�9�-���QE57�Ɨ�9	����[�r�R���5�v�2�HdZ�M-�����:9]#�N��4E��c�.����9�
]���٢�g� ���s���g��f�s��-ֱ��̧K��m��Sr��jɨ`Sr���wɘbS��̉ɈdSr��I�xfS��́y��`NSr��Y��gF�J��9�"��aJ��9]$��aJ~�9�]b�ӕ�2s:�f?�+yi��h�`NSr���%���7㮏�?w����9��ٟ��W�}x��d8�+�t��K���/��K!�T?]��K�ӥ&�d�.���{���K�ӥ6��=]�K����A/���Aό�C�3$���G�Iϊ�\���I�UIϪ�\�����B�j�\/�Y/6׋}֋��b_�.׋}֋��b��bs��g��\/�Y/6׋}֋��b��bs��g��\/�Y/.׋{֋�����r��������r��g�Ŀ�o�����p���x��|��\���ngw����s��{���H��>�c�y��C^����ӌ�/�O���}�o�i��/����Ì�xx���M�շ�O������?��_ӿ��TV'+�z{y���~���/��%ʽ�8���x�a����������������ǫ��<������������-��������@Qb�x�xs��}�����kk���f���D��(�ʺ�>x�&��N�͡��W�>VVhB�}�֛ۇ���p��5�|}uw�?�]}�:��>O��}eM��-k�\�:|������+��JӔ���{|�W������=M�B(��;������-�Wf�^�ik:��5�%?��y1*�s�+G��v��b����+k�\C�r�)�3�Y���~˵��,ˍn�Xn���r�\���<:a��M7/�ir����_�7w�N��>�[?i����E�p����7�������t���o%�'�ғ��u�No���alGw�Me�0Vv��WCj�k�i��c�a�<���p�m6\��$Kr��H��B��3�_��]�r�!������o����~�}��7�^��ҳ�I/���It���J0o�=�,T��U����nNoL�_��}�l����*mbpb:w��1�}��Vm�c%ߌ4�R֊*N��Y]u��KC���=]nC�-�SݼxS�Ow���K*�\sd��޷/L��>��D�3���u!�*��ƍ&6�mS���@������ZU�P�N�u�&���kr�_��X�]r�m����+�>��;]�\��x�Iw7M}~�m�I������3���C���kzr����Z����.v.��4�I��u���6�3���v�.����V�S����j���:���S�n��Չ#tf2B�>�hB񃵦uO������o^��k��M��Pț�B޾>��7��7���x/��o�v�w����>_8�ɻ�������u�Ӈi�w��6:W�����h�U�w�v���n|t3�[��xj�+;;�r/5�Ҟ���K�S��}���W��-_K��+����&:�T{=݇L���W����|�ZWud�X�Cն���m��a��h�z`-�������|̫�ԯ�I�;�g���˜���^��'�uj�Ou1/�r)��zi���Z-�{j�r��'�v���F������.��^u�ԙ�F��o�>��o��?&u�~H_P���a������C�4��s~���������_�þ��������}�����h��������տ��OI�W�?�f������������'a��qA�tY�$�����H�(���~���}���q���?�p�F'�2~�.�uj�ү�O�;�z���Û�3��^*��X̵+�>���կє6[�tU�7����jf�{p������ظ����G�t9jL��.'��g�v��q��r΋�v��y�i�زU2��}�*.���al�X�f�t���}gS���Vq�f��}>��bu�\��5�J��#g�*���-�%;~�)� �g��A+����j���XfXi/n�.�P�5 ��I�W0���`Y0+x�a �=fZ}]�-@�u���ü����S'�.)V�մ+�~���\~��E�� '^�2/�-d�3�ͩW�_�蛫�x��Y1\Ӳuw,��ݶ~�E���^��X�瓕�׉ʳ����bu{_������Pk/(Vh��^d��Ƃyۥ��u�`�V%s��y�Ud�F�J�Y�b�5+��M�� v�1����zC[�σ����:�6�����G|�b�o.S���U�R��>��ka q����&�F�%E@��������8�1��H�U��N6�J8�ֵm�z]��,�����q��!+����ۂ��X���FSv�3_�Y��Y�fy����)x�T�j���Xө/��Y������t^����L�T��l(�z1
^�BOmn�̞�8�=r�lIYIi��6��m`��s�Mȝ�j��ٹJ�&\�q�0����pv�quPӸ��5m>z[�˦1+U���w�x�ܲ�텸V��,a'�¶���X�����5��x�JmYm9-^}��V���z����u��&�;(�m��e�!��:/Ur=��+e�;C�^�U��9(�N�������m˼�0ؕ��^(U�Ԃ�D}�R�.��6o��7hぷoK�[��8�۬T��
�i�f�
��\�]��ػv�	�O��~:]�Q?��B3x^(,���B� ����ȶ-�2V#���`�����q^h���vs�]tt4�=�.�]�.�]�Ev8�P�<4t�u��T�ez���_����>@�ڙA�Y��3s��5�s^�Z�F�v:o-ŵ��om}`�/.�4xyq����a�6��:�wݹ���+vs���q�����W�e�����h�Z�h���Q��8΋qk�`�C7"k��Iͭ�����2�y��Z���bu�e����[o���y������Zg��n��\�-�u�g��Y1n���?z�������jgG[�-�Y���>/V�oٝ��J��f���XiD��!^���8�!v԰O�O(��y�b���	�z�[wt�q	^2\�w�j_�V��N�O(���X���������!k�����(�k}e>�":i?�T�]�d��g�Ŋ6��� 0G�;�8˖�}�7���ݼ��y�_�eˊ-�-jf�L�R�=���\��߭M5��.�����41�<�cb�b�slM}A���B)�g�����Z�x9px>]��l�.e]g�g��L����T���Ŕ�R��#�Ηp�񆃸Ÿs��8��קo>���3`G/\tX��kѱo�����;w�/�U���vֱ�+w�}�����7�?�e���q���??\}L�����;��������O~~zH5��׫_�PK   W�dW)<�4I � /   images/3f348383-912a-4adc-88a3-03f2846ee105.png <@ÿ�PNG

   IHDR  I  *   �]   sRGB ���   DeXIfMM *    �i            �       �      I�      *    :��  @ IDATx��i�m[v׷��Ͻ�����W�����U��-vr0 ӈ G H@$���1BH|��H�P��D��H�$D#��l�\ئ���]�^����~����9�^g����q1��{�9���͚k�u��Y��/?���g����{~۷���w�ӿ�������?��������bkut~�\�.g[ �W[��-V��������b{wwqqq��X����۫����[}�>�|��������G]<��s�Gydq~vm���\,w����b�{�Xm-����|�\^�-��,���ŵ�k������������b{g��8]-���V�R�b����b�\b<ΓS^�&|���� ۠�'d#G8	�d�G;I!�~�����w{{{���}@��������xuvz������e��0�#�(r�-O,��������_��899Y����&��b�+�Y��/��֍'��B��Ν;��G�_�+'�����][���;�彿܋�g����-
N����^��"y�n]�o�/��GGG�M(_���zXQ��I(�d�B����vzV-�K����,���o�NO��h�<���%Ɩ��z��-���L� E��N����۷՝_m>���'>O��'W>��.���ٹ���n�j�<D�&���6��W�?=Y���+W�,�R?;;M�߻wg	o��^���Z���n��"��+�b%�v����w�F/<�4B��n�?�9���>�PO>�/>2��Q�����h�9���+�.l���aG�߉¸�}y����92쏽=&�uv<0K��N�����8�W7}m���b[���:�?�������:~-t���WDW���;���7��łaB���	壣3P���d;Q��3��ߡ�.R%\���+!�0d��-�7�T����/�����k�v��۲�������6��R�����t���ߗ�K� �m�+���6��#�X�a�ko�2�G��e�t��2q�kms�m�"Ϣ<����ޞ�Kڛ��"[��+۴b9�V}�͏�x��]��"�Gf0ԇ�Y��C���[�ı�L����ła�p;����bqvq��^���Z\ta�/>���u����~\|	#���.�L��G~xh� ���ڄb�Ʃ���;X����� ��o���g�������L�/K��F\('i��ps��1n·nz���Ư�������h>�s^QV��wVo�?��ͽ�+����c��[?��g�/{zq����5h��$�w�'[G����}f��Z ��SG���I΍����NF�m���߭As�u�~����0�0���l��8#.�W������إ��܇��L�������l5z��ú:t�n�h5�U	fof���U��TG�|�Ĳ�'ˢ�ƨF�����	���qr����)����9�8=[�bLwv�qY������L
��P��F�����Y���.r;�}ᢻ:_o��cP��6-���m-
N�.�T6���QC
��	=���܍,ۤU?����ei�3�#��;���\�=�/E���b�ē��w�W�l@W��D�n��vy'��Ҹ��,u��f�1�2���&�_L��>�ϔÃ�B����Fd�ۇ�e7��|u/z���u�C9ueJ;O�;���day�~�T��t�����+ֶ�)�t%��|Ǧ9�u����Ą��-�J߳���ڳ��1��IwA�:?;@�_e���[��g�'���G��S����,
��k�V��C��nFWg玓��*n`M�Ib	#Ԣ����ԍy�e�}v,�o��.��o}��N�T�@RX^Y����v>�Z-uq;�O����kR.6l��e�bSpq�<��r���lurt�<>=�l���KU��/�����'+�S���z�+}b{b]j�^����GiI<ʫ���G���E.R�<�2mP��Ɗqh�a����K��"��a��~Zq�U��L}�*mS��苈���C:�����ƥ����"�B���O�܅�}�b7�yϝ�69>��?�n��'3)V�`�?�����Y0n���]^���$��vw����O����yA��5��q�:�M;[��]���,�h3�)��儵���`�:f�<ٗl��]��g�gt t^-��n\�[��o�������s������So�k������u���b.|�F�a"���~��Z4��0y����k��|'
�_z��w���~��-n<�CϞ���o����w����lY�\��v�v��G��\:�����k�S�9`]D�d�qbdӲ�Jwy�֭l��x��k���:�:4 ��]pUb'�H��W/NO�9��`�s	.��Ce,�0	�_�V�\�с�̼�k�SOel�);0����c�wA��gu�M8�$�9�X��tQ����f�A{=!��|d]��|uUo+��I���ly���䕰�����W ����p��|��#/&��dл'=��<��S'Y�B�=�l��)��z� I�[F���lcb���Y�IF����
�.�H�ݲr��o��A�1'-):��[�a�c�l�P9n�G��� ǉ>���f0�?��g.8�I���0�'mG�#ò��Ǐ�_���ú�&Oqv�&'D ԫᚬb(W�����q���j�۰��G� ˅H�Q���Sx�/�+l^�S�l�B��N��9e:ܻ��e���
c��c,91��o�ǵ�p����P^ㄋ%���М-��O�c�h/N(A^D�I�Zl�M��g�1�H��5�����,2l�_�29��q<�O�	=5+�.�sr%H;�G��
�!w�FBx��6�eێ�:�l�x����L]T�3��_u2�談W1ދ?.����y���ݹ�fI��6'>�����Prq�âxrt'}i,���_��_�@�~� �N&�Q9��f�����v� Ɇ��.���4̝��$!3��G�#��x����� �='+_>��\�;�V�v9y�6�S�.U��"_~&�ԍ�13?������ȃu�D��O����~~ʾ�Y\W���L7*�P��
�G�1� ��v�;B�zl�V�;W;��+�S��e�������
���2�/�	�Qc��W��~e�^�_�R�ġ�#�Z9]C���]��z\<Xqggɉ�����ŷ��=[���w�ݿw��7V��|�7��z�-�A�q�z�!$�S~�����i�m3.o�������.훥���7l�������_��?z��{/�x�������-N�^�`�m6H,�\]r���s)���<�>[�ւ﬒����nwa�;��lO��>�\1��{����wJ�вkw�w笸�vq�n�8�ʐC�)�t��:	u�i�ౌAJ8'�b�iZ݌9'�L(J��6�^pN���?|G�G����QB���3(�&N>�k�U��	N���&ٝ�����y��^��b���u�v�W���)�?���������Eh���!�*&P�&�/b�*W�LM@I��4��������,�����b��n5��ڭ�m�����[[��2̕�m���$lu�/�����#�-y�3S�Cx��	E����gn��3b���g�[�.֞����D�K6� p�����=�C�؝����I�z�ٰC�'[���2��4aLy�ݱ�y�B�Fہa��� ��e6a^�N2l'~�%|O��`Xl)��ӱO�iJ]�G��~'1%\�y��<��*����E�+�Z�y���<�n8����l���M[!��f]Ӂ�l�F!n�sE\�eOb��fb���O2���ٹF9����č A��}��ؤ��l��~P��Ic{&_79�pNߪsӌf��������e���v�U����)}/�S�h#��m7^����؛括���$$ks�	���+?R6f�@��w�N�LU����)y�[M�|{1�g̝]����plޅ�gGs���|��qC���n}�8v<cJ��|�Ы��	�OhrڥO$��4B����M�u8��G���Q�z�YaJ�6�r�l;Ɖm�������=��\!������Q�>q�>e��
|��.v�j����������Żl�-o��=׮�{����_����������������O�7�Yn�H�p:o�y}^���m��&r�.�w~�W�/�]���������O.n�>�8޿�-�k�Wn�`ﻵE/��$r�~�U��){����W�d����L�̬u��q��՛��n<���Y�r��bko�En5ݿ�Q���?���Nv��c��	�W�{�A�� !B0q�V�~6x��A�r�M"�����<�T8^"gq�H�er�yX�F�靼�����I�L:I^U�y�٤n�Nh����5�<.���q �X�M��]0��#��7R�0U��,zSB��e�I�k0��̘�
�V0� @&�8k1g@4>��2���6��Q�������ok�A�7O�f�V�Jo��FNRN����������|�^�H�-�M=Pǧ���h�D��P�(X���.>v�g������sԎ���/��O��b/W�N)�d"����\2���ܩ�%ʣ+��c�r�{��+�F~,+s�Ѳk�Ӌ� ������ܱA'�����D���H.(���al�t��S�*W�q4]fD����j2lcK.��{�==c\6�ʋ�2�,[i��ihO�* �O,R�ȗ�E��8�زYD��J&��-3C4�\9�#��A�H�B'-�+��g'�S*i�6֮����5����C�����S�ٻ�!g�g��%$5.��y�4|�\�m:��6������#$��7�j���5�ѫ����������qZ��+N�q�f2�����$�e�?c�����4�,��W�Ȩ��A�p�'�Wz$H�'y�>`�`;��	xXRB_���t:�0nlqN1wYѕgؚ�:L�� ��9��f���of�*��qs��'���zE'p*/��n==!5q��p��`31��~����UB��6�>��5?^���A���mX�/�*��6#���Ƣƈ��3.���y����1���9�g�,^��g����r�7���|��/�E^����t��9��wJ0/O3���[�yÄ?��a�����Y=���l�_�;���-n-'W[�|�bq��560<�ѝ���8�{e�$��w���r$wo�{�`��q�G�����������������{��9=�����+[����4�3������ �Yp�`�8'b��I˝���|.ƣ�&mo{�y�R}Do�h��q�<��u좐4�f��pr�V����AI^��@MW�A�Xs+�ܶ��G�T-���%�s�+U5Ɉ������6n� �a�&�;If�+P���P�.`�`:�H����"zrc9x{�Vpi��^�����9s�+~�;Q�~�>��`�+���L��e����I:Z����i���Q�t򇥢Q�/Dۗ��-��IR����7�¢`h=C�,�>	y��v�aM�:9!��E)|�/6'�'s�Z��e�Z�t	�ru��h(���ĳ�{�
-<(h�*��@h�[-!��mx�E� �@�5U";��Q4z�x@�	�����`��| 91�j_�� � �;=�p��PS�ȧ(V��e�;ƨ3�T/o��*�XNP�O�e�q���ehkJ�"Џ�Ͻp���iFg�g�8��x<Â:Qj��#|�ciD��Ϊ#ѹr��"����\�]Wg��)=ȈDA�'��c^D�w�_U���(�5��$����O!��6������ͤL'��\@�@	��)=�(->G�RʿL0�����b�����:e��$	\B$tĕ����25���^�B���]a�G<s�?H9�@cS�9՛Rz�k�C'��bu`���4��C�Wf�)�R��V�U.��� 5���[!�:c��ј������{,JF�~&�����t�8i
�?�q��"M��>��,��@`��,�֞�e����Z^�z5�mn����V���;q��`0��a�|�ʯ�����ŗn�^��ח���}��Ï,~=xجg�;�/��no|s�^��nzk]�j��ָ�y���Y�íwjz�w^ۿ~����O-�>�8;8dWuy�����~��z~-�b��~�k=�Ƀ�u�x�7�e����+0������g�������������W���l�J׮�_���b�����o������j���Gw�?X<ó��3��M?xĭ�ɘ�I������p���
��Lo���1Q��N
#�-��z��ԥz�R���Ddx�� �T"���=p�_�s���v����M��8�Eo�2S3����:��'74�35ڑb���I��P>:�Nf��X��<ƑŝF=���4��[����B��I�\d������0��Z.:��-�)R'��g���NR_�;�D��%��4�;T�w�Ղ
֩\NIM-�	��I-4��5;|?�K�)yzs��W`�1�P`��K�uI��� +�ʚ�_�R�d<c7�e���Iɗ�-�@2kNڀ&|�q0��B6� ��)�Z,��VT㡞]I�$����E���W�nB�u�H�z��;$7<��,��FR<�u�Y�1Nr��������@8��EHu�(����(�)�3������<\&�� %�Ϙa���WnN�����NW�E�06�r0�R����F���G~\��A�;I|�B��̕���kH�?T2j�;_Y��t�֓
aSl��+��j�9�֧��G�
��ǜ�7��-�Tw��g,n\��HI&�J���Ãg�hL2���d���s�Āi������d�K���{|����lzN98�sI<P��/I�>P�V���s�K�z��L�AP70*Q�@Y���9�R�B��Ixd�V�|�PT�����l�$.� �r��]�o�v��_�f�e6w�Z"�6�Q����R&M�3�zw!����^���r״í��㛱�6h�		W���O��P���0���6���o_�`n��]=�ڭ�ѽ�o������i��O�̛|u��l��MPu`p6ۛ�&��Wk��7�[�;?��>���+�������!?����_���|~�x�$Mǜ�����bwq�|�HO����_�~�ŏ���o��|�#�����k\ ,~�Ѥ���_����`�����ϗ�������k���/<�;o�����>�-~4�:���7�7nN�N$NX��K�K/]����6�N�֟�0��F�����p��_�I��)9-���<�J�Ev�\�~�Z�)�@���r&1�����A`�u�Q�Z�8{3z�c�+�"�+��(��^M��ȟ��t���Y4�x "�	m�N�	c��|�VI4�o�6%ޙ('Ɏ�zX���^�����.޴���J�$��_�Z�K�熞�y�I��Q;Ϻ��S�U
p���(�>a)�p��Q���>�ɕ,�B���bP
�J����G=�s��=^9=��z� 
�nH��郚�1P�����|�� ��D�p�u�d�W�>�Ԫ_��5�5���A�[/� ig�*���,�Q4́�p�c�tc���NO숒�E���eMM��[C�n�hk:��ꈳ�a�o�f��7u���STዦ,�k{�1��g��Ƌ���T){�ey��V�ff�G|p^�iW]�S��%����Fc�%޽��ך��xE�/`��,:��!wz�u���"��(����|XG�ڂ=���Mb��m�"�c=5s|�5�s�7θ��i(gϧ�Ì|m`��&��0T��Og:���ϋA.a��H�٪�(��)�W[�;�F`	�}N��7�N\�J7f�yJ��B%&��C�)�(�y��ۥ�.x�IEW����QI�f|�kn˼���v^��Գ	Yq���K�􁖺^PfU�x�����ǩ6h�X�x��ƈl������M�	��J��͌\�G<��2��3 �e�I�(�-��>�1���N��Q7y��+Wxh)Zͅ��[&#��^��X��������!�o|�ٗ����X�0��sU��9\��s<��u��7]�k��׹��4�7�9}�>��w~�_^����[��3~G�c�Y/�\=�5:s��-��q�vvg��c���>y��;_���~��������}�S�.=�ՂͿ��|2?�+���_��j�w���/����_��?���������;G��L��A�^!x�%+	:�\h���p�d ���Te�ئR`g)GX���p�!�e<P��m3� �j#(�RG�F.l��=�V���'����w���n���3a��Vy�ryf�8� +&_�2R�����$O'd�J�$ ���(\�^2O��.��?�w1��S#�|h���n3���P�L=�;	��������<��N��	���8@J�uN�9���S��99H;p7G@�i�
5W�p>�|9Y�+ܦ{Y�+�鸑X�� _����T�J���Ƶ����32�I�ۨ������ �,�eb���GD&�0�G%�̓_�%�9�����O�uW�~��<���3����j���1l�߁�v�lo��b����@�Ej���X"@?�~�������ǅ�FBt��R��Y^p�-D#rʜB��{(�&���G\E��o-x����b�L���:�Mb���`����*��DO�5 �u�>�|1�:	LRZ��{|5���<i3^��C[|����ȯ�>���#�`Qc�A��tH�0�Q���>��f��M��6c��˅�*��^FCP�F�
��/"�u}�"�k����XW!u�b�=pD���m�.��ӼZd��w|�+�b V�7=�$e���޺���%��ϖ�� ��pH�-��8��A�^.�n^0�o�S�v��/8)2\�	�s΍8A�|ǋ���[w,��y���<��z�/naC����_ء�'��ǫ;�W{�{7x�@��1��1��M�f]L{���l[�E�<O������&|�.�ג�s�xdu��`y�e�)^76ܴsӋh��7T�ʄ�{[�w���+g7�Y��̏��������o������@�+���u����S�����˟�ħ?��>����w��s<��K��6bPȠv��u����_�>�$kg:N�dDR�h��*(pۄL|�G`�6˃��LX3k��g�)�1�a�f���>0-	���i�oGc�D��L\r��܆��J����"�,T
)�5T�m�ѶffC�7`=�;���G�[��^{���؈�N�ۉ���VqF�`����������6��)?�&un%���YL�Y{�Q�}���kˠ�n}£j�#��6�j���e�m�c�m���v��v���ğ�噺��KO�P��j
-P�i�k�Y�+j��>&.P��<&z#�	�K���f�C�)e!��3%�BS��n��@\}�J�a����=�_��Ȁ­+�y$��~��sxD9[<�AċoKOB
�c-jȿeQ����ֹ8i��!�����|&]�a���9�Y�5��3.nx�Sg�;²|	��Qp�S|�?K~]���F���p�B��pο�:_��X;+�RN�X��N׽�ϣ���q�'�:HZ�zS/���5rZ�?��o�*�ƭݛ�������~��w�'�R���G�5{���`� rSf� ��y�PD���Z��%|df�T@��>�r�`#.��ڙ8&��].��'B.ns� �G���x�w�X�w/.���v_8�������'�_{�����{���/����Ͽz��_;^-oq�����3v�_���Ý��#^:�	����ِ���������q�9m͐�-rU��Pw"|�>���ZGjyR��s7ۄ�ۭ�FҜf^�vSƼݶ�kW�F�\a��}E�`�5@W�������w=������~�����?���_�]�z��BMs!]nE$貧L����������~��#���O>���^>��8��o��� [	��Dl��c��u��\��Ӡe��K��e��:|�J�7n㤗�8q�6-���1���wb>HB���}�rɪ��f����;�<H�%�|��96_�&��k@8���(����2��c��>	��a�RL�Ǳ}�gǎ>�ڒ@rx�	j��U�?�!����l����T��91��u�ɐ��|/��|rh��)o���[�݄[/=&��+���g�+k��{2]����h^'�J�I����R�߀�{ֿ"KC�/
Xӆo�zp�_<mY���uV�sX���F���������m�vM�]���J*K�m�|�P��
��)e�U�s7Ǎ�+`a(�hp���.��)�B8���:5b������چ5�q�>�t��Q��:>���iH�*���ѯ�Z"ef^�	cA���ى���U�6�v��<���[{��
�J�f��aB��;G,��a�x�CfN!rs�ټ�俞��Kk
����`<���2�x�/��p�dmuғr�5���8/e��~��ԙ�(�%���H�ps'/ƝO�Q�o�+�S,���R8�EGɜ�F��
�q��P-�h^ڌ"[�]�>X<q�������������WW�8�u���ѿ��w��o}����w}�ß��߾��x���� ��?�}|�8�u��g^�y�kϾ���^x�?|��W����ڷ�;??�>�_�a^>yp[���Cn���k���٣9י�ٱ|��aɸ"i���rׅ���>�w;m^;d��`��4Ks�]�����.��w���$�@w��"�O��1����x��q?���/vo���w\Y���ş����G��<���9�VX!o��8��>���ſ��?���G���o��?��K�/�}������Xz(/M��5	�[$C9F��d���-6g-����A�4�k0�����@��T��X6��K:*�4�O`��9� O!I.@�"��2c��)��E�'4��i����6�sp+�rb�EX�������֛��yW����6Vh�\}9gMV�Zh�M*�Kydd��>�'MdY��u���vW^���L8�7S��nS�y=��"���ڄܴo��oȗ��O�f<��}I�����%�%�,k�L.vfT��=`�LϚ�v�ЅX^�A:Ÿ��b�ļ,�S�7w����D�؝�k���}����vep�7G%��m��N�b�""�d2�U}��S�t��֏{o1�g6 [��v�\�m{�z[Q�a ��Z�'T!���t99Ǵ{�������CU�|������>qh׏wX���e���R*U�7�>���ЌÖq���
i�O���b��uFbjȟ�Kd!��S�+Ⰳ��:'�ga�0��g�xN�?�ܝ�f#�a���2���w��o��_��~`�[q=]�h0}��ۧzM�5���@�#��(&ct�a0J�\@�����m�6����eO��:e�٤\����������s����/�o~��7������;w��[��7o��w|�������o~������a�l��S��Ͽ���g������W^��go���_�}�;�Nηn#����.��o�c��x�ǋ&y(�l�'�IG3`���&FaN+ͼ����y�����چ�)��7�+ZD^2ã���ɣ�����Ϸ����݋�[�m��_��['�/��?����iS����I�.�?��~�����y�mOݻ}�w^{q����_gP�X�)��w0�=`�*� C3�f�yo��!�κ�D&�Zj�wzri1��/��(�[J(|i���&����w*��|��1��F�/QvP�ŃЪ7eW+�fREK�J��%�zh�#V}xwltj�}"۞�+�l�%��!��÷��y�'���v˳i�t�M�6�V�W��b�-�'}�~m�):�.��_�u�%��-�����;�LWP��0�	6�"�æK|XJb�|$2w�xiJ��xD=(|%4�G�e2��L������So�%(eU�¸W��_��̦����E�AHQ�ntx�H���s�`�E[�����д�3���FҜ�Jr�3R�|<�A\�:����[2ɍ�P���Ґ�DEL�Ѳ�Ү�_E~�L�sB��^�_=��%��l�M%�	����j�2:�~8�
(,sBK-X�;}���af��R��cm ¡u�<�~6H|鼮�NA��������k�kW9p�4��yzD fZ�<a���MQv �uB��|MS%M�s��u��&g�f�˩�{L2��y����7����A�_�&���*���q�чvI/Z(~�(ϫ�U�%�s�ps��XW,v���;V;�_�����~�m��W����ӟ����˨� �f���M���ަ��<���O>�S�o��ԋ�?��_{�5��E�:�,d���p�ju�rO��Ѭe��⿵�)2�^]V���yi��S���q6in�������~^��L�Ư�}T ���$r�x��������?�����,�7��@�[�M�M#Z����c�o����?�m}��w���������O,� w~y��r_���&����l�*�vT�Yg q	"�	F��舨�OZ�a�V2Ŭ�L@z���I,Ac��j�uQm�cp �����.*����e�<��8��d�q�C�GT�XeP῜<a���I��a��Ͷ������X�h  ͫ)y�u #嬁r�1|,T�\��V}%��9j�JR�H�hI]��a�i"���S��1(�uU�љ���R]�N[��fa��RA{6�ZWͮ=��T�y{PF����z��p@u�}`w���� *Ǎ:6��#t�>�!�hn1�e^�b$U��7��f;�E.߭b�i�[��F4�����H;j�'�)���c���R���ڏ�vy��Ms(5)�ܮR&t~�z&�{�yV�Kp�"�|b�щ֓|(��(����R�������fs)w!��n�2~8=̤��B�Y���h6'�Ci�_
%����#�����T�;��Tr���e�R�f�C����s��6̃��Y�k3��S�{��<�LgTB�n�ԧ��/���:1g�1N��O/�5��E3eWa�VJp�4���y���ݵM��΋ ����*��c.�A�|��[.PԻ����<|�s�N��}�y{��á�5�{�1֗w^z���+?�{���������/��!֌>��@�|�����!������������g?�xy�=s�����y�<������$�<��uȸX<�Qſy�&���NZ�y����_/�;^��@���.��"hy�=�쳸�K�����~�w���}�۟Q�VH7��6`����e��i�s���?����?��g��������������,,W<'���UE� �hl)ꠐё��ơCh�)S1��@׃^��0��K،v��k�Ueٻ�����(¼3A!�k���>R勼p�;htc!R��)	TД�E|\���ׂ��r �E=�.R�kJ5��õ���[�����e�tiv�@Y��FA~Z����N���Ԟ���ʸ��4��hGI����!�d	j�5L+�薉����v�yb��z���7�?�N�247���O�Zٲ^��4��W��a˂����h��B�	��%�z&R�S�/���B�-v�uf��x���%ԉ�!?����?/W\'d��#N�{���|+[@b�����P0���'���+A��j���O�z����2NQ����s��;���$��4�X��T~E)L��FU�4�7�Sح5N�i�9����$T~P 4��w�{fHd���C/p]�h�)޸�|&+GRK�r����$�2~��2y��f,�^nN���Ώs(±�s��f�1�,i2� �ɽ{�;wn����{�:�?�xr���q��}�(��UX|�Кi@��lx�/�6��ɻ>r���
H���Y�d��̟��<�o �^�V��F�i��ig�R��
�u�OyM�e�u�%�}ō|���PrŦh��=��L�%�������+���g~�/��~���c9��������ˊ�K?��/���g��uz��'�K�{�ݾ�_Ǹ[+��=�l�bo�>�(�L����^�#�y���w���_/��>���͑�Kaz�7lא[�s��[;���o����"o�k�ms#ۨV��M��9�?������Y�&�w|����n��g�N��c�R`�S��S>�Ģ�rL&iO.��B.����5����ц���33C�5g�yϞ*���Æ�נ,�X|�\�����<�	C�T�'���1�OV;a,39p1�Kj��h���k:�U��m�z�u�9��=}P�1�㸗�>*,�C<�<FT�ǏZ٩	��ǆ���:���3����w��+�u�ޜP��|ӯ���r�>��������V>�g���ZSt�������Y<�����u;�z@cQ���|���V-�µh#��U�*ۧ�m0Շ����*���;��q�b���N��r�L�s�U�:bV���ݴ��y��ֳ��.��,`?��[�7���$T ���ᔀR�(�`9��'�P<�$�M��4�,��u)Gn��)���4;
��/��뀉ڑ����o����� ��,����NVr���"m5&F��?޼-�$��;k̕ɗ��9?M�g?��Y�P6K�>��b����Jf6�o����+������<Ǐ��?h+/��ﲠ ����α0�q�ؑo��Hf!�QMe@w{��|�G'����¸Ƒ{��7E(g�R��;x怃�w=y���������������t�Z��g��nk�9^�~�[�����G��駟y��_�a��e����:�;7������FiJ��[��W���I��)'���_��H���p���|��vzs��÷,?����Nރ�����tmh��ۮMC���������'>�#O���|���]��{���1ƻ��A�.�\,�;9���Cdbe�k�i�=&`/7�T�w9��8	�1��������ղkS���5J�JtT�/��#�w��L�Y�g2*��y�6/z�">�D����B�q�u���q@�A^�P@�P���i�1��I�Y�������������+p��߬�it��n�v��L9�4��C��y�_�D��9Ak'�����V����OJ�j���:5��֩yH����s���C� ����Df�j2_�Խ@�d�C��-Ӫ�]d�c.���%c0�:#4���5u�pm+.���V
�����,Y�@t��;�e��ծG�)��~ԧ˃�q��������Z�F�[K}�,[���A}�ա�c�7�1,F#d������s��U���$��/��D6�k<|���_���!�F����n#&���?��6O[����8���r�:Y�zUn}���<>9�k�LT޼�ް�I�"��ϗ����|�U��Ы3��Abwe�o�֮)?������g
k�P�.o��}�R����4�������]_U�eC��6���_�o���3�K������:/�o�\�1n��7R=�?>{�\R��и��ʟ�zlq�������~ׇ����Tگ���'?��/����x��_{�S�w��S7O��o,O����Y��W�=�n�W��J5�,�|��s�g���H>�����Ӄ����ژZ!��\�O�]���W�]�����7�d�F���/E_�=LH�5�8��ݶ����_y��/}����Ç��m��ݣ��ސ�1�W���6��N�$@峑3f�jz��k��'�.�[��D����V��%ȣ nh��ǁ�p@�	G��c(B��ĕ^�'��i������"���Zh`�	"_O�Ɣ��ՠ�O�mmJL�"��t8�:�݄2&hpKxs0�����?�mȉj��5>��2�CO��Z��qa�}��d�.�˯�hfk5���f�j�В�2���a0�<x��7��l�]x�s;i�lt�:G嘖��ُ��u%IgW�k<� P�Ħ�;ZsZd4�*ZJ�Jl�F�����-�	��c�W6�/<�6P�,
(�m���X�F�T�"�fr���  @߿/��9qr��P��-p2h~��p~u)V��w����~��_,�4j�ʑ��;ſ[7��xH����9��!  @ IDAT�.���bذI�mQ�� O���&5�Ų�i�.Z��������o�b	�XGM�m�N�+b"T����VP�n��s00�?���~�y��D����-�������lHʶ��q7�Qi8!��Ϟ}u�FYz��?C���h0e����<Ī|�/2�)��ҩ�$��ए��7����R.*���V��j���B�ߓl����}�&o@�_�w~�xz~���O]����?�鿸���DY��I}ߐ��v�"���v������ϟ��ދ[Gy�3�ܾO�G��o�gJ��e�zIV�~3u�\�<o����375|�_7�[�2���x�?m��t�NW/�y�ի��m�~�p�+�ٓ�m�ȳ��37��<=�f���o�v�-�=�o�}��?x��՝��w��e�T.���TV������cp���J}��J��q��e����u��e�0�,��gjT`�j ��i0�N��	�$p�ɟ���:��$�SW�'\����f�!ĉ����� �UN�^
%unP5�=�3u����8r���bS��_�	�*��Vc�r? �D�a?غf�;�GR�My���_qi�U�'(�nr�j���~���O�l�j���u�͵6�3���3~������Ք� ��x�<��X�,�5����-{C��|
O����\��_���"���:��� ������&#A�bU;R=(��U�Mɻ,�Y�������~ ����0��d�4ؖQ"�,z�o�.���w�Z_�S���R�f�!�
����[lAf+�Gԭ�=�a#��rh�8�R���Z�=���D�>��\<a<�A���l3�"�Ri��Gm]��K:e��µ�1F����1R'�e\$��W)��G�ch]�(t&p""'��X5��N�FB�:��T��#���ډ(ZDc��u�'툩%������xU�N�^cU���M�p�>�ɧٷe�e����^�Н�p���s^4Ed�����b��~��&����?����?��o�	������������/<��Ͽtr����O~�_�����Iw>�ݽ����F�G��r����\{�}ؿ)�#�\!���w��_���W �N�Ň���7�n��8	����q,�~�c���_�z��;�ۺ���K�-�\1aD�_���J�H.��"p��zbU����Bov�(BXںғ�z��f6��T��c����|w<�p *ĉ��o����P�ϻ��.wv���!�>�`q��o߭W�.�v�5'ɤ&��Pto��GX!�)�|���O����f�h���iU�:�U�?�2\�2h���uHV���<�T��b$C�F�m6��Ϸvt��{��o9Ifc��o�'���7(*�O�xN�"��}p�y��oV_qԗkY{�\h�Y��vq������T�u	ܛŵ?ף��ރ�vM~KB��W��6I��]o$����ș��N�,Ր��^N��i֮���U�S�>ii�q]N`��Z�󬽧�]����D�;�4�R��}�j;IC�̡����=�&~�^E�m:��)�
F��E�4�-�H/�vX��/|$�t��'L�F~)�d������bcP�>g���̸r�W����x��~y���V�����K'Uy���<s�����Om��fY=�=�m:9=JdF����b��v�_�v!.����_�p>%ы?���͏��Ι���Q'w�&�ǟu�>���dg[�ԅ�a͹���������ū�!�q�:���W�+j�#��Nn�_{�����;�.6���W�v�'<+|�˔��'�|����?�}�����L)�QO��&�Yۀ�}�;�5M��8M��o��sw����ć>��M�B�K�����c�lr�ռ�c���x��fm�+�����λ���ͳi�>Ǳ,�mǓ�X]�Г�K�Y�n��p_��oD��9�,�f���B�83�i�~�v�w�?|l�[S�%NA�p(�(t�M���ۚ�R���	�����z�FƘ��~�e�ʷ崊���B�ֺNm�8b)���o`�x@�.�,���L�W��n39�A��;��Y�F1F1�������ۑqdD踕U��)}��Nm?�.}��+�@�^/��6x֢�����#��:`<#�N�OW��N�[�	��pa������_��`�ߩ6ɰ�3�� �w�+�<`c�X(��#R�2�1Iw��3i�7K O���3_�
@ED����+�,%�P�S�EOF���+�YNB�e+9�	���E�h���,X��.�2��q%_u9�CE����҉�')��|���.���
"2$����VH|���89�����'8�n`9坏��R��j�~х�������'-��E��
���х�nN�X�����b�ȑfU����"9/�/�	K�`ۂT_�K���H��As�!� �H�,3�r�5�4?���]+aw ��>��&	"��|~��?3�h��鹹��<�J��)���A
o�]|���g�ZW��?�S�0�R��rϠ��[����"*�OQx�|�	J����s����59��<�׬�|#��I�Rf�_���s�~����<j׶񿳨K�[̿��:z�}���^�7vO=�����/-���������-��������~��e�^�*�v����0��M�yÃ𐯷��Ƌ�?��>�ܿ��������_n��w�;r{�����y�b��l3������\Ƽl�f�i�]���C��%�ka�O���r�{x|���s�����lօ��ʿNaַ�?�k/��dV�W�*AE�z�\�8a��g��=�K�A�9du�˰ۢG �\��,�~�ơ�J��K�/�I��I�z_p�U?��� 9X��4�ZG.3n�u|µ��F;���#W���2�#�G2�MQ!�Ⰶ�A�3aW���(�Lra���ɴ�e�~�ȝߣ���!�%������M�3��.�Z�uC$�s���lzS�*B��J��֟�=2��t�Q"*�*i�`�ؼ��ʊ�n�ӕ0���lI��X�rW�\�slY��K y��b���R���2�+J(���`h�5�j�#K�*
!�M�����|�1͢������й��b�7	d�Vj}UE;���s�8��h )�~�W���=N� KqL�08�����\~������G���KDx�!��˘@�Z�*/��DP,�� h�ch�R��Z�8wS�K�r����{�A��S�SSٚ��+bz<�aعE���ꋭm�Y��[���J�{�2�
�Ȯ_7�ܴ=,�����g��C+������s��H�)�-D/�4iw��QEjx䏓%���ñH�d��7x!V���n��&Eok�И��!<�B6���t��V��7#��A�����|%�"�|-?���M>Fj�՜�e�r�����*��F���׾�q����+���������Z>~�
���ѭ�W��;��#�!""۪���6�״_�q��';��\�p���c�,�p�E�2'������m�۬�c��ȗל��s�r6��LMk��pl������?�}����L�򛈣��Wޱ���ox���<���7s�*0��B��cj�������?��/��2~��f6����ɡV+�,I�0�'�JT�ֲT�dru�ɨ5�P��ep\
k�N8E'3*YVP��@�����d��d��۶Q��,"��?r��\Eg>��`#�����!K��|�>�n���rUt��i��̍�o�\��h��	G���e�,����c{�m4��xN��&R��NU��n��]ec��.�D[x��hC���Y�.��@�p���r�Md�2-�|�m!8e2�#��@�����W�A�x����n�2 {�א�@*="��onKfzq"߂��̮���Z����Fw<��ǇU+"��J��6��mk�6-�೥}u��|��eŀ�wY��&���~��t��&9�t���u����� p����=�1��	�5Ry���UӋrG+��v�Ac��M��j��Ff7���KL�=e�24��)G��ɶ|𣙶i#%"/�Ish'�J���a$t�{���-I�a(R0�5�C'�/T�(��n��)�%�4��GX�|X4����ۆ�T�r��aj�ƦۄOm������Lx�u�̲>��a�FOע&�Um���p��ٰ�ٗ�ʼ����{��������rş�ɻ��s\[�'���z���^9|���ʸw�O� ��s񢞅����������<r����>ד�.��{����1���7�/�j���y��;���0�-��ݾi���c��sX�t޼���s�������$1G0��-7�O��sP~������/?���5q�>"�a�|���y�|�����>�"��Ƶp.��)_	V2L`b���Q`�z��@թ��߯|��B�����xmU3��#$6�d��I�<��慧��>��I�����A^�p���m�������� ��_���`��U��,�T� 3�+���y��v���p2يG�M�-YD�mRfRь�M0�98��́/s'��0g��	�Z�Bh�C��8���`�?�	t�aa_1{)��
*�
���S�Wqa�����1/�X�t�:ox�d�.���8�o'Q⓵����$t+�G�MAڋ��~q���Qr��"�|T])Q�?�G��\�Rf��<J&Њ.��uTuaRq�=J>���x	د��q]�D�0��!+L�}T�n�_�k���3�څ�B<��[���A}��RG�ԁ�ȝ.
(���Gz���.��24"RE ߩ�*�a�F���	r�Y
��$��I�!`3=�̊F�!j ��V�p�s-3�D��rVO��U-r�Y�8�g�1����ԅ�8�Ln��Wq	�%�V����-p�5���V�Nms�׼����l���0J�
g�O3��r����� ͘Y�+\Qe���L�lh��y�_:�vQݤ���	��YT�=x:��n�w���KC����Պ���-�;�ó��;O�� �3/�(9Q%_֋��'f�7n�M�8]���r����7�/xK�s��������K��!�,�4������w޴C�ķ��m�ֲ��y�v.�4�W��n�����p_q��<>����;~v��_�=:��i���/}�`�eY5����L�9�t��4s���~�)��CNTXPv'�I�+�0���x���]r��1�2u�f}��5�'B�1ڥul�y(ۖ4dD��[�c�D�C@H�j݂�M(М1!��RΖg�ǫk�]���?�6�2}�	�'Y�8�(L��Ŕs	:�P�,�i���CtJ��ko�ֽr}өl�Vm
�ԅ'I�W�T�F�t�h��	��"�+�����($��Frir�*��$T�$/�Ś�U���������']�ֲK���^��6xM�U�зh˖��@)��3�i�"�����bR�mQ6����M�8qhOr�`؆w����\i�,���$ ꛴^30-��q�5u��a�Ie��+"l����/�����.fc�M�u�M�(�InqS�̙���vr�\��h�m��<��}��u%�@SՉCf"�&\��5F��P��Z�5SX�4v��
��<G)���t��`�L��Hsɫb���3H[_�qs���5���m�e�E/�*��Z�`:@��D-�Ac&��I9.g�`��h<�ɵB|O��7���PrJ*�������r�p/�|�{��`��`y�>}�SO=ۿ.��c����;���>�5m�M3ǱL�'��"�n���3�� k��p��ȓ��� �������	��7�m�&���:o�9�f�c��@�C����>��<ø�ǋo�,�=���|�K_��O|�We�g.���s�_��h�;�ܼ���k�^���1`��D�qq�
������fm(o&�.��1A~	��s`��a�U/?\�9�%ZRV_m���P
/�"��u�@�u�q�%6��!\�j(����>C����6��9��O!��6���|�C��G��2�'l���״�4_ U�0���Eg1�X�A��������I'͆I��f�Io�������6)hE�M�n��q��%v�!�h�6U^��r;?�F����!���!iR:����y58��������i����9��ڐ93��s޳r�4�V�t�kC�����	��G�1@J�
� X��8K�uE���#]Nz�h��'���k%���T\Mu��|�*b�#7�E�����Ǘ�'�!�.o[:զ�k���`y�՟(�������K���5���o=+/?���Wi]��|E��''4ܾ0��g�ڎ��|�w�	�6�ͺp�ݼ��m�_������*���6�B�X�S?'x�|8��k\�r�����Gov\�w9�Z��'yk�9��yy�Nٜf�������+�˽CN�8A��꾧�WO�]��m#
s^s��������pf����y}5<i;�i�����B�\�lWX���[T�f^q��:����{pp����_x���觛�\ʹ�-t^o؜ֲ���e�/�V�Ͻ����[/�~kq����e���e���_~�4i�2Ȁ!l�Nt��+��1��3�y�=f�!�0�u��XN�P"�@�Y��>���܊��ރQ�խ:pJC6���U4�#_�O`�
6�U{�������h�f:�LcҙF3��3Wl��R����z��B ��ņF��/���PLX�
/����A����Ǐѳ�N��7ZǍD�;�&^]�6)Wй̔g��f���i~���@b��X�<p�^����v���������Fl.O=0��o��A�I}����
�4���JIM#��%èN:\�ȈB�%���ê�%�6��c4�9��p�v}"A��[�C��x���m���<�7��ǳx��69��ƃG�� !o���z�T�����}kS���n�H�Ql�}�W�\���LU"��F��5kF��l��	�L3^T�:�c��a�d��^UZ�J3%��ʶ҉�����@�T7��}��D��]L1�����h��r��� 7E>�]�zߒw�8�|xx��Z�T<�Ľ� l��N
�.7μް�p��.w}��s����{�w�O���8u������[Yq�^�[Um9k�ʀ�?���7銚��*��۸w�ͩ���? ��7���nʳ��Y\y��xqõ�~곟�#�Y���J�b��f�i��]����_��Wn����'޲x��x��?��HU��M&^�pH�mG�*�ܰ�; � P&x���6�y�ds�Z:~��DDwMʬ�!�vϡR��*.����4́�3�^f G=�C��j���\w\�_�)�'OY�(�>m?Y����g]�ħ��[X_; ~�^�ϔ!/���.����~�!�9��O�����sG�$0)�:�B��|�V��$�˧x-���Z����Sﲴ��*����0��?�s��>1����o^�t�Q�n��ěûM؜��K��@�4��(O���j(�,����p�����;����6a���=�d���<#��Qvэ����f/hx]��0t�[�i�M��ؕ��N^�#7~Kfr���W�R`n��l�ޏ�:-cYݽ�ҍ�h\���g�����cJi~�Ǻ��5�<��/�2.��~��9Ǜ��׺)�Zt�9����_��;�ě�����-T �Q��ߴ�W0��;���ǔ�x�f���-?�ы<��=�l�>=����W����{��ut��KiƤ�n3oxl��m�n����˷{���o���\�u�����#_y�����H_/��E�mC��>�o�����N츛(��aq����K/-��9�So��/������[U�����f{�7�����x�"]����?��r�}��c����..xh�`���,?TΏT�A�T����npM��h'��{��뷺�^��z��Yf��y9�(D�x-�H�^>(ldU#�X�#0�$�\��y�%s��4�ș �IedN� ���t.5}$_�+.��(g���ށ�p��,em��,)���oD�(>eԚAm���W�\�����<�-���'�N�S��A�q�S��T����P�}��� � $mT4��,8�i7�&V���Os˟��g�Ha+�'D>07�c���h�4c0������i�&t{���xS=q�E�����O�Gy�����>��'����������)X|?�q���~���S�R0�����G�|\�>� "��>�MLO1��>f0ħ��?�p'�j�E�*�u>�W������.�n���B0¥�tJ�9�+&�� ���QşzK"ݥ2X��W�5el�x]:i�}5h'�wy���9<|�y�qֹp���e[O~j��W�m�g^ބ��,O����� ��0�m�~��2|���1�y��Wb;��fd�9o����2�I16wv�x������j���;[�߻�۞}���%��ɮ�sf5^��o�Y_c���t��O�����}d���}������X�����+̜�vyS��������i�����}S����F�!ӧֱ�w���V��v��ʹ�O/��[��\�\}�;����G��?���y�	l����Rb�;����?��OW;߿���~���s��ϐ=�" %$N��(ʗ��:����H>�-wgw��X��a���2����h��@&ܲKz9��$J%���S4���6K�;_!�tIY֊y�(�����m,-�6�mw�C�1��DY�Ph�.$p��&�`�ɘ]���r�l�O]j�@�+��Y�2%���Ueh=��rOɥ��̙2��>qP6���C����Y5�s�{����c�lT|�كO[�	s*��o��|�А�h�ɖ)�f0ۣ�P�C�Y���ۋ��˴*JP�{6�'K(4M`Xv٪�k�_�5c�Ot�c.�ȹ�Dn/d#Qu�����xF�y��M���̻�yú�'�BW1�ms>�o�N���\�E�w�<N��s��g��\�N�ٶ	��d�f}��Yn^���)0��Թ�#'[�X!M4�ܰ�c<���yd�M9�	�&�ڦ}�Z]Y|��,E�C��Sx�s<�O��wT=-<r3��s��1�����}��W�u����>��-?�8�M\���|�z��g�����䑷��=P���O��C���+R�m��]����i�2&OӼ�a����C�Wí[��붇��~�&l��<6sq�s�zqzqλz������.�7�;'�_��->��S��~Ӈ�_����o������s�/B���M��)p޶Y/��������Gϼ��v���o:;�V_�������b'�|Y�J�$������ૼf4@ް�mr��y��~v�N��0K�H넜�c��tz�и�iS��E�j_9r�:��*�2���7.bs�QI60PdĂH%^�`�.�M��FQ�$��԰ʵ[���}���\7�r	<�KѼ���<ڷ��;�ww����ƞ�՚'!�yv����1b�,baXLN�����^X����qblLb1H�-	�uk�Q�z�����/��w�>�~�{owKH8��v�v�N�:�}I�����P���D"(Q���	��tp5�кfg���bk��E'c�&%��B�Y��,�UgeîQ��Y׌���$ǃe�kO�K�H�ں:3#��7L�1�M��˴9r�u(J`^ɠ��d,��E�x�"���*bI�,äv��-��*;�G��G��{%jr�)�QK��Wg6�m�����7	+P03BЙ ��|PJ��X���,�����:Y�Wy
͸�{uCm���Z#�t4/(����I�GA�
�ƪ0pњc��.�\g��W�\���e���]�y�VE�/�&���|��򔫪fY�����W���{X4��0Xi��Dh�N~�+a�U��r=�������@U@�k�͢�pkkk���Ԭ_�+�|�Mo6�o�>�������w����C�	��ua2��D=�d�c0������g�_6\X�����\�yK����-�6����_2e-#Y}��Wҋ_�jޙ>�<a�����<2��j��n�n�vw�}Q�Q_���7m������>����zus�����������O~������d,�>.��T ��U���7��|�G>��x�ɏj>��Gu�Ov̲���%�xN��5��W�(>�7 +Lq�'�z�]�����k��\��l	�+���0~�JQ�(�x\�8:���ʪ�s ���f��G/PM���:��1b�1����E�iǵD���QV4U���3)'��Ir�O�NS�qa��2J=J�sF�|03-�Gt��}�zY���:;$��S��Lw�O �\$��'�/�Iݕ��0n�=x*�@B�4�㘮2�8Bʍ8���`e��0���|a��@
p!
qD�C@����3�.S�M��9�O;�y/PJ�)�K��v�b�4
�Q|\:U)qVRq�������K�q����_)I�G�S��RF�*�t�cϒ����5*ֵC��yĠ��S�tZ�I��?�uܮ��ze�����]Ǫ䓢�y<����O�����{	�W�?53����5W�^o�_��<������G����^�U>���o慧�����G?��_�����w�q��$����v�ov�3���m����_��8�SF慣������t�_ӜT����>ed��eIS�Ù��fz����m�m�;������r�L�,M5�vЬ|�V�/���G��;�w��U���?Z�~���o}�7�&8J4^�:�Y�Ǐ<���m�ᛦN���ǦW_����'n�6������p�����
 ��:8zz��_�KS�v����x�8Uє��������N �d<��� �=�}nW�z$�n��� ⥑��S?n��^�T�-~�L�,:hq 9:�7��9%Q#\�ǳ�RH�+�Х��1$T?]��A���\^nlQbzP��/�ŢtbDRތ����蕜�����p����_�-��K�����oW+n�&$i�V~j���<�9Y3���ԛ���X��W�A�6�#�����^�Ծb�_����cފ%X�<V�2���/�xCL��������O *'�x*��W�)�Qo�X��r`�,#eF�X2���/f���D8.?��p��C�E:_�f��w�����3��*�� g�E|�v�տ�R$������j�E��4������,z�
i"�$<����逻����<��)!���{�+�#�h��$eG)�XF4���ۉ�x�U1����%k�ގb3J�X]�� �GI$�ʒ���!���C���-t�p\;>���h\*Ü�D�RE�p%�E�T������;������e�I.�Z?4��b3�|a���(�����^��j
����:�=x����Zb��y$���]�}z�����\����Wۭ��|Ngo�1�P7h�s��x�K�����B�?��h:+O�^�kxP���_��._^����|�+������ؙj���k͍�s<�����]�;���&ق�s�H~����eL�O��O��e	ϲ��Ϥ���3g���%M����x�`o	��~���b����?j��Zo_�%_��g�ٹ/}�������O��/�گ��'�^�sR�:�JT�z���^����+?�3��?��N�37�>ojny���N��Gm��Xk�O�Қ1I'.n�zP�jY�3?'Z�L	 >�qF8������R�:Tp�W��n���N�${q�C��!�<�� TpC2?��T/�8X0뭞��
�]։�{��]�tK�e��q�:N�q��ϸ�sR��.���d�Ƕ�UM�&�����	�&IVy,�OJ�nA�8��l]E��"=-�\WtP��:P���"�2/�`qϬ�e��`=E���rNwmQ0'�q�:v���'�1qǇ�D��N�,�&ˏ�ulR���I�^~���ɯ��Ev�m��PX�����ۢZ��7�S"7�s���c���ɏ�0_�J���3lLd�(����[�_1��N��Z�� �	�BK��U>n�G��BwR�vG�O>�\�~�K677����G�"C�L��V<�/:Z��&�E�C?���W���^p�6��.6/�l8��z�Bqa�����S��z*=�o2�|�O�Qy��䷫?�}����ֺ����O�������i��[���ۃՖ�s��u/{�}�+^ڼ��~��z���h�y��}�_�/x���|���O�u���N-��㎏Q)m͝�xm��͵�<�_�~�>��#�ƿ^�򒗟����^���׸���G�nn�G;����=E���YK8�/�8$�rKK�az�NN�9c�U��+��W3^��0�B�+���D琧H�A\�|�e�H/=y{� ��#j�	��64��꙳�6�x��^�]ia�H�O:�N����̃K�������Ș�CgQ�Ԡ����`���qH�S,��C҅nt�,���w�qz`
=�����N�<";���/����ZTڀ���S������˧?I&�3Zd�W��#����d{*�Sk�N�`ٞ%6RI�C�;!�I]����D��|�d��v��m��m��W첆�x�&	-}��(��}*�D!+3Y'M"	;b�$v<a�$�q�O�E�<�E�k���V�"(仢�s9kPٿ��X��_Q ��W���?kRɯxתN�#4Z�C�jZf9����~�yE�Rsxw˸X��B��-�����e�AL�b�3@���;q��e^�t�^�cK9���+;J�l]��3���S�U��?莁�'�C���wΟZl�ڽ�����p栝�6�s��`m�n�h~�����������K��?��~�Z5�}ȓU���ě�/���S?���~�֭o�ʯ��W\�9m.�i��O4￲sx�t���f��1:�w��໾����R{��%_��εn	S,�ꦸ��կ����E{RHں<a�}&n�\�΢Ĩ�E��=`�7�o0é����ħ���߿����o^���k�.�3����f��?�̕>�ۿ��ff�/��n��/l��E/�)������.��Ω�Ņٵ��3��;{����/-6���V�T3s�|��w�����,�]h�YA��u<k��"D����9��.�y���vN҉�r`g���z\����bYd��'��ֽ�8w`ja�I1�p��:^���p50PU�76n�Y:ľ�*ˤ�U�r���N���?^�:�p;-�I�3e��|�&�� �i:8�#����@5M�rl['���z�����$~����/��r����y�W�:��ɻ(m_xN�eL~�#��3I�|��9"_�u�m<�}��-_r	"��$I�vY��XE�ɇGҍyl򵐞�X�{�S�G���	8uy�հ����/b��#�6L�x����Q]�?������SԩJ�d��u�a�#��N{J��~�hf��n
?�EE�q6�W,:K��XnD)ٲ�~��=��:	������ַ���|��	!}5�2XAb��D$�PQ7��刏�3�6W��h�>���˹ͼ�N�|��us0�!��v������/|�w|�7�����o}�����Ï�&,�	I�o�)9^@![>���������m/��~�}��{���/~��Ⲟ��p_��#o>v�V�?{��	�,��x�m~nf������{ɑ�����O�*/[�G����,i��3�螳�IS�G����J<��<q���୼���}�lk��=�-���~�R��{�n�������t�v�f��>�\~��fv���__�e{���r�讞93��9�N��w���6��έ�KW.7g^�|��Ï=}yp�����_�\���7j��`C���ď���$*F�ɇkόA4aTX��1���@/��.Wh"���,�<qt!��C$��ϻI(HO`�Ip���N;GJ�F�k��b���Cv���e'���CeJ��ֳ�Gѓf+���Q�1�]V�*SH+�m��Կز��8���Q�Dg�Т��ߎ�WN�N���q�$����I����/��"e�(_ݧ
�K:�U~���1	nfi��eB�xI�AA'��v��|���_�!9���"&�2?]�?�-;uQ?�_�&|���AT<�7&��# �3�t'�.K����#�O��dP�����$]!�"=X�]R�[��ˤ|�@���$yS�n�L���JL�,��Q�K��x���q���$]W:�kh��E�J=���W���F5c���L��s�<�����Z[)��1�? ��!������R��6���������)ʺ#���]|Q0�K�}-�8�����Y�KlD\8���n�l.?�h33��,��so��������W��5������?������}���o���꫾�O����s��VU�"M�W0����w���?~�k�~�ɿ�p�ܗ<�Y���U���T�S�;>��fg�ls��o��Y� |>���ы�������W��[�&j�����!�K?��íq�t�c��8^�;�G�$}�[�4���������h�ۇr�!�ՙZ/�8�FC6{�jy��<��iM���r
�gx���������F�x��u�b{jf8z����D��w��ln�6O>s��c���ի|n{�nRs�����v�P�m��;l~�O͎�<[3�r�ٺz���������s��
.�v���?n e���Up�H ��n�L�g�z�Z�Ȇ!��)�(Vg���$�5$��B�z?!������R�T�.$te�E�FgΝo�vې��й��ђ�j!�zv�����=(RM��a��Rٯ,��]`��ѭ�c`��>Q�N�^~F�r��J��X���"��V���T~���L�}r���ԟ:u��I�$���U���c�T5o''�����,�_��?q2�q����e%�$�゗<R�W�!x4W?��܆̷����$uY��*�ٔ68ce��B���O���'�~��n����#��
�g��S�|�Ȇ���vU�'�WH)���{�=M�zȑT��LP����|4M[km��&T�]��b�4U�w((�Py��#?ȇ�]���/߄��}���B-��S�� ��"����	4Nʬz�@���.;C�k���q`�#��$��/p�Z�Gڹ��v���yni���8s���C�ac�f;���Íf����V������o�������l��_��G�������G^���z�+_���_8w��K����>�c.=���ٳg�777���x�������>��_�f������}σ/Y��}��M7��F��77x�k�\{ȑ�C��E6;F��i^���֟�������f�G{L���w�I�5�Nw�U�.��B��WdN�T^���$}{�/<|����n���s �ျ�r���L��(��j��P������E, vo<1��e��{Os�ӣ{Ξn�/�4V����+W.5�[|0�`tkg���M��n6Y,�.WצG3���pf��F���������U��K5 ��T�<1Z�Y2�ET��e���H�h`Ν4`uW'Ɠ�(�ޛGx�%�W2��$��mT��Yr�YW=|=�;I��(ޛ�{��ťv���I:L{'):7!)����WJ�)r^�0F7���§��\EQ�-2Q�!�U��K>�ˀ�p�t ��Ǘ��6mRxOS�/�,��u:�3>��$x�e�xX,�㢄+ӥ�")i�ʔ�ڵ���5})�a	�;�R�%vV��.�ʎ����I�8�g�dʲ��隶�?�=5��O�X�O�&$��I(���"aL~�	1�&�tKXQ�pxL�5�O�����w�\��&��`��5�s�g�"��l#�%��,�v36?X7�pr�x̾= L��1;�l4�@JS�*�����iu�M)�l`�}��f���r������g�NN�����p2�gU�LT�k��O�$���0Cr^TJɇ���3��$)N��y�V;_��&B	����?s�t���$�©Ņf��[�;��ܾq��y��]kfX(-�q��y�}����C�yG��o����k�?������oݾ}������'f�'_��?>3�yfv������w7X�;ܿcko�nޜ}/3���Ϝ��λ��Y�m 9@ƿa�ͩ���NӼ��k���n��J3\>��4�<5h��<�_n�pߩ�|��|�_��m��`��  @ IDAT�>�@�e*��w(/.uY�N➸'��O�OV�pwwG_�Վ�j����P�-2i��n�Fs���h�i�g۫�;��s�:o�<��+�+�\j>zu���ǯ�gO-4s8���m΀�3���a}����K�[�����t��-��S�v�6wq1vZs,$��m��]���8���W?d���g�%��@T}�Ikz����qcQ�y�(?��gyYg8��ʖZH����2@����nN�?��'F�_��\qG_���<eI#�B�#���Ǖ��uz��L]�I˯�k>��L���<��|�[��p���8y��:���&�Is�|�F���M�I�|��r�5�d�4E�����k�Iu�N�lj�1�L(�u�C��\�mTg���Ft��~RF���c��G��1~�E��2�W�Y��'�:_��|�~2�4�Oa�O��,��V=�Nɣ��g^~J����`.����u(��Ch�4Ņ�/��:������K=��?'b��e�{���?
�%F��V��j)>����"�,�4�
�ő��Q[d�-���#A��$��4/L��4�3Wn4��sO��|��{[���ڸ�Q���ы�ۻ^����{����������o�֕'���ǟ|���o�瑧wf�{�K#��{��X�M�����l^\8s~4=�ୠ������Fs����C�?�\۞j���5�L�����V^pI=ϝ;מ�K�KPUD'<��lx*K��E�t�E��;��q�f\Ó�q�����!/�jfؽ��n��#2Z �O���L�6��u�n�%�9^���Mr�l�]:�!��f�7�skhj�4�P	S�ay}(zF��Q���!�0�E����|���:(����Bcl�� ^$�t\��6S0Tq�O�(2�U@pSYF���lb�	����*�q�+���G��S�i"#]��WKR1�U��T�QR�$p�)d�t� �o7 Dv�6 �\_����Vp��慉Y;#���A_A���y��q-D�̓,��U'?�G~��gI噐#���+�BU��l�R~D�i���b`�y��Zr?�P�E+z��.	�S焑��t�;�pT��ʋ�SZ7���E"e*��N~>揝TO��V>�dĆi�Z)<NvM'z-���Y��0K���W;XT�<��F`?
�E�D�4I��Yg�3}D���-�R�g[�PC�����t�~4fC��c��. e�j}�ȦQIT�R�����v�z\�2KA�;�y���J- CDl�QD���`q�����h�����6��O=�)��fp��?��h��vuT}8��:��֣"
�wM����U��zۖ��^E�� >��E>�
�t1�A6�f:4�x��h|5B���C>v��g���%6,vvn!g�o�i�Ȼ�g�Sw.7���c��W�7����~�+�W~��[ׯ̬|⩙U6+|~�;%;��z^zqzv453�m��;Az��^���As�k�SW�xv}�.�R��f�N{����|7u_s��p�裏�z��+ z�?�]u�b���	��N�|��`*N)�,�3G�e��<a�y��K�pz�-JV�l��Đ
f�R+��r��I��mzp8��8�,�ts�E&�D>-�-Cv��#���Dk߄RO��;�`c�K��<M��
e�������;}���1�_h\V�8	/�2��QMJ�kt�н���R>C�4�#!7VFF<6�X�	W�'��#l�q`�O�K�.UH�d,Y��|V�$=�R���V��I_�GB���n�2P@T���I~�ķ��IxY����d��u8�o�Iܓ�T��ğ�'˕w����(��Uy�V��?�NY����d��u��LZ��i���4�14fPY�"��ۇ���Fj�oUX�l�R��L6,e���Y�qW��1����ʐ���\�xZ���B]|2�r�anf�3B��
�[��m��j��}�1�^��ݝ� �Q5�S�΢Rի��`BK�X	߱
u�[��������"�C�� /hW�p�A8łD�m&�����셻�W)߸���3`�te�&��G�˧�|�t��=ּ��'���y�޻�s�gGs����a�?�7Y����˫v6x�͵uv�6Fj8��K[�Wy]�5�6N�����:��_�'�ϋ19:3��}��_��Φ�Ӣ�Dc�|�L�u���'�4uZ��2�r��Yej�m�e����h_ ^���@Դ^ �:J�lQ�M�-��!�޾-�hE��i���ם\����g
2����~,0��r����_B9�öɩ����%,c㪎T%�'^�AL\A�Y.j/�Գ�S։�ð��"����������hڔ~� B�Q=}V�|]!ښ&S�$�_����4�]j�:J���ǆ��AdZ�OƉ�y|c\�h��&y$��ϸ.Sz�v/����Q��������n�
��D��(0��h?ܻ�?e�/>	/t�?u8�l�����<������Gd$}�¯C��'N�o�|�%n�(NX�u�ғ��x�O��W$,��5��@HEF�I��$�$^�/��k��`�w���讘G�7q���r-�D��o�c�6Ak	�enaZG����8�w���	/��zˑv2�ݛ��pv~����6�/h�4e�j!��k'YBeZti�!�����W��s'���E+F����}����u�D�{�� �{���Î@��N@�����նٹv�ٙ4�����l�.�nv~vi�?y�j�.5KYY䩹�S��e��X��Y>������m�8���n���{������
���v�ö���ʎdYY�C��ԍ���jV丸T[�T_�	��`u:�kx�S�Z4���d�Kt���隦Ng�x$<�?�jR�8��;G��:q;�+b�vϝP���pd�q5跳8�^ (�-�t�� i��\� O݈V�C�A@��Ad/?�@�K_6���(�3N,)��ĝ��|�6ኻ2*�pUK^�X	HO��2.�I;h=V(X=}�z��D����caC�A:�&��89&����Ie�#�3N�:����q�	˸�0��+�3N�:����q�W���[��[e^�`�I�:o�'ٿ�-�U�R�)Y�qQ�ɺdyƉS�w2>7a��5���D�����'�d|n�2��$L��W�v�xu��[l���׳�\�?��'�*a�*S+M:�Yό�:e"mU�HZ���O�>.��}*y�܌��k$�O5iW+$n��UU>�u�nH�\���f��Ü[]i/���z.�0�t��U�A$��J���Xe�Α'�#
:��l� �t4��Ƽ*!��0�C����0�(s�y�����pN�Y��jW��E���~���с!��6�b��M^��Ԉ'�O��1����a�	�cbc����#޵$�3,2�g�v��9�?�e�`���hw�-VQ�!/)Эd�y2g����yo�>+,N��T���X��f+v�(�,P�M�h꼬��^��$C8'����'��y��p{g��f�Gv��%ƽ@�-jlR��lJ�zssM���j��{PY"��e�P����x��@�����)����U�!_�'����O��8K���K�ɸ���>�M+N=��`�*� Xo kmoӂǵ��=��VJT�J�K���B
|K�:�pU�d�K��KsY.p{��B�q2�G�:��;�Tq�d���qE�d�g,`���W�t�d�����{�Ь�ߐV9?iar�&/�O�c�b&
w2��>�K�E^:t�U"J�֐>=�p�O�=E����`����1E]���;O�&~�*����d,S�N���Q��h��9���E�$�I<���g��cqf��y)&p�iW[ó��`(VH�J}��&�c&��D�u榄1�Vv��Ę&��z�1>d:�ޭ��2�d����ǻ��v��A�OϷ�g�s��w��	���)\�9����g��
���f�:xw�YY�yBb�
�@W��_�Pd�'阳Զ�>K.4��d�(��as��NOO�VVϵ��s����^��!�g���S~zȉsD���S݆�;�v��ف��<�:��u�ZɝK��Cfl�=38D�B�v5�A�^���Q�2���5�希Z\�����`�eZy��|@��n�H��%�L�<2LA8�^���e������;�T�r���E.&!0����W�<4+m�6��8+.C���0�wmeUs9��1�*sT��%BҎ���8j$1d2Z7b���t|�ڥ"ia�Jgx掋e�>X-m��t�x��8��~��*濚�s˗�>X~����O�?��� ��>&�0�J�zN}��Y�{�>uD>E��OV��?Y�G_%ܮo����?����A9�B����X��}�#�7�.{�v�?����uz���?6�����D_)�D�1�j����/9�T��(*�]:H<�����򻺇����������Iz|m�����މ�祰��`^�i�B;���ޘ�sYK� �6���Yv�ۼPO�9�M*��?�G]]Hvm��9��+�6��j�c,`|����_�d�'��}2:���eI��v8�=7����v����g�w�����|�{p7/�<�Gr�x%����cWL>-ORf�?=7+ц�W3� d;�Y�'�9�=bq���v�8��y��M�-���]I#^0�])^�'.�
��i�c�����<i�K��ʞ-Լ���ϔ�!_�u+�Z�6�[��{��)��d)�G�����l2��X��#o��0}_"���${�v���q�u]2)�K�=M�~�4h`I3�Yje� �+V��;��*���g0�y52� �D��xL����^~8V�>]���)z�N�@�hh���ue����Pd��_2^�Xp	qz;�j ��������ֿ#�Sؿ�Q'?m�y�2��:y���Ika�*h��l�������I��:��W�����4i��?e��L���!��M�SnƟ���u���ʧ���E�o���!�;��D�d�3�S׿�-��~�+0.ߓ3��&}��A��Q:�P�?��c3꜋�n�$���:�p��\'���/zו,�	�������8�^`�ᤌ<�0�!�rI"�1���x��c�A	�q�9G�]�V:��0�F��2T9�,���{e��5q��i3�#�@��.�o�!�Vm%�$�{{�l��
�'���q�v��r�y�/j�7�5׮]�ml����é��ª�����a�����Sc�I�1�5��p�n�ۗ;�Ӯ��_�0 O�q���$=Ѭ�u���;��;Y�#��g�o֥N'��k�:��	W<�2�2��`
��ϔ|m��HҌ�s#yp���}N�s�=�j�_��5�c��Z�h�_r,T�/��]��i� oۈ�݂Z˕a^��o���o�lE����%3��K��D����w����O��ꬮ\H�5?7v"�Ǆ�N'je�3�r��t�|
�~���2�t�$}��8�3�����U��}@K�"6^�W��:�|*.�j����+iؗw�o��r���}����t�3�_*������g�W|3Yˬ�Y��N̴��U~�.���_ŝ#]*��0�j�U����ߏ-��N�h�/�DT<8 ��;JXzO���<�Y �EvD���!���Ȕ��K�%��9�,��!��aN��տ���}�;���T0V���!o�V_�+1ʻ��j}ڋᇧ˰�`ȧp٭�~�&�z��l�m6�W϶�y�g��G������[�q�z�[���ƴ��΍�����z�����Ӈ�Y�����Jl,�=9+�^��z�ss�����F���0SG�g,[(�xi���x���ĝ�����q�g,Z�/ye��l��Zx���҄<d�4����&w�؛���lwx�Pc?g����o�T	���6�yj�X�j@|���;辷��x;��z/Rڜ^�K�hUEb�)1ȕ��z�{ǀ����UK!,e��c� $�
���3Uux�)������zġ���Q�8�������>Hj��;9�<cn�?9}ф�s�!$�b���i��h$s���+!&O��`j�kVK���Sq#�76��rg���k����<����(U١�|	9	�4�z��*#�n�dWAe�c	�&�L��.�q�J��Ϥ�'÷Y��@Jt!Y�x�u?1�Є>�#]�940������,��;��E~�(v;hk�Y�_S�㣊��h�Ѧ{�tc������5�B��,������o�8L�*0!���A3�ʁƮB��;vad*U{��Xb*�a"���o�]l5�� V���'�
W��|N���}��� �i�f���>]޲���Aԟ�<�u좢F�a\��r��FU���Q�qh<��*p��qmO�����|��~�H��� ������{��}G"֞�*��s���mv����C��91#� ?4A (rı�"^>�e�Eu����s�����"����,2�FG���n�!���R2�v˜3[v�xĞ6C�֟f�l�rF�C$����e����C��<�|wY(M7��%w�~����`��i�)n���{��uO�,t��g��}
���>P���4;C�Ц�nY��
�)n�i8�n	3�ޱ��#n�1�
F#p |��c��O�I�٬od��쯺�?d,�B]��(y~�5?����gyQ���M#i����}Y�rJ����-��穪B���G;L1�j�Q�3�vZ]gw��cF���_ܡ8KE"�T��Kg7�R��\�W��$�9�з����z<�,��|-l$'��H�Ś+n�IE"�\��ę@/_��]}�<m���
���$���iJ�/	4Q�J�� ���Ġ�oɇl�����O�TK��?�*r(�{@d���a:B$�	Ծ�z�H�)��Q`�+u�\:V
�o~� I^�'݁*����,��X;��hVU=�1�� ��«,6s��!2�Ȳ���&f]�#�O�c�.*CV��?��#.pשé���
{ZҘ��C)*<���%B�Z��K^"�B�f&E^���$1Q�	2���{�)��LJT��K.#�ൠ��]�vb�*W�CM�1��2�5�����|R"�՗N�$�w��L�����,��'yM�?្��'RL!{��kӦ���v�@�mY��2O�_ԉ�Oc`��O5Z����w�I��?�f��A8�z��YO4Q�	�����Jˢ��oFȑz�H zfe��(��/�����n���7rO�.���O��gù�э���ԭ���3i�n����ܙ��[�pa�E��|�9ھ���gY��?�ZeN�R����$y
�u*m!}KP	=:CB�O���e*WZu�.WY�O�B�K�5l]fĉ���e��|����ܸ��O�_��8h�b ��X��8<��m4��� 6Ƹ۬N��[lR���MWn�p]�����jI�_�L������zı��Zu�e!-4�n���jP����\�d{��x�@J���	���h�Z\�Eeh�U=%�Ž|0<6��23��LR4�vT�v"Y[�FZZ)B�����M�%�|�u�Q{j�R�ȋ�eu�ЕE����y�~ʆ���VH����9wI�z|p�21����NFϰ7WW�0p�M{�)����S@�
-�n2��������T�W�30�Dg��Sٔb��u6WI�/�W2��<k�-�D���IG���h!����N^���!�c��mJ}u���-�c��M1�^�;�< hb)��������TL�.ͥ��%;����c��K�5D�1�I6��{���z�^3��ڹ��	�ڒ�\!x�X��R����L�,K�*�6@��R������'y^z>��,�p�}Ɠ��pR�K�c�`^�45	}�x�;;�Bq���]�+�6���1����Uc�放Y�������Q�U���#p�t+%�g6�z�,�[ȭ��V�'�"�3G26fdV`=8��;�T�g�x��<8��(��������V��6Ѩ�j��;37j.������͵����/������:�S���*ǹ��-�C���J?�a6�}�P,���sRPi�e�Z��]�8vt��Wf���)-<�w��&�I��|�DGy%ͧS>/0��S{���+3�6��㐴���bP����(:���L0�0c�T� %�~�S"#�\U�i�i$��g�|�����(+��N^�q�JR�+�����;�H��(�+�rJ���r��:��ǁy'���qAs��ջ?t��4*��?�|�Hx��D�搮X\��� ~��%���!��ab"n�dMQ�v
�h�R�ԧSC2
b�7Kц|��>�$��B&�v��C��b��Z�f�Ji׍�$��m^tw/���2԰Ӆ:T��v�zJ��G�|��*��$I����VL�w� 1��N�'y��9��n�E�2D9]�ɲ1��Q���3S������a����]4��ʽ��BҠ�%=��l�%m��2����⩝Y]Jxӈ2.,ʒ���;���r6%ma��;�J�l��26 ����u�"\{���D݄��P�o�]7���%T9Hy��T��,!�c��B��xUQW���pk�:-��F�S�N�� Y�j9�w��rF����.ʗ7�[��K6����[轘V�����\�*MTZ�K1�rQ:m={72V���	m�:[B ����+2_b˗��8�����b]��p�V#�o^mg�څin����~����Y��L�N�n4���g��+��.�<�{������y|zi�uѦ6K9_sp�0�8��܀~�W !;�P�6�~����K��?\�W�a[�@����`��� ��|���hO*K�䟼�q�g^q�L���8J��.�M���$������h��|HS���@OZ�>�I5.�uC[��q�A�q�� ���8Mt����l�� �ؠx�����]P��nD��O�|�	�#$��/	,�T�����ǆ��X�H]4\ƴRYs�R�� ���V3�f�k��+�bd�چf.�����ۿ�5�vИf�p4YJ�[��5K>*Ã| ���5#��ɾHd��;_{��F"�$1 ���	T��N����B\
�:~'�2�m7N+(x�)�I/�v�G���Y�.I#x�׵�S���>��]��#��X�H3��c�$���K4!_������b!�D��,Ҋu'�av`�JH�1L��[���r��U0������K*�%�2,�^
^^xkT��� Diş[O��t�de�QWc�#Ɯ,g�Tq��D��zJ�����ʉ¸a�~X��z,��<*��5N���.+Ck�yX���P��*�PL�X�cr��̃�i�M:���܂�3m�ߨ�E�8/PO�v�'����HJU,��"�%oh�Z�O�(������	�X�����Z��\��*�Sp$�\����|��`���2)Ӎ��Xf�E4)?V���-��>�� ��߷ '݀���`ꊢ�+ɷh������K���+-{L<�?�-�
����v��xʏ[mw�m�ۭ�k����h��v��nn eoks4�c�����`{k����ns���S�:����In�Ȇ�3qD�D��ޝme1��qw�����UR���Xe�'�d|RY�~�>.�<k�5�I2DW���7�
�S ��G;��?:�Jj�lF�-�^aw�ӳ���0偘O�޷=f�bA\�gGzqA���|��=E�8�%�:�-�z�V��0:�����H�����f4�$D0G�J��Z\۞ ����$���K�V*��gpH�"�vn�}t�F�9Q'̦�3��c�C���t4U����y�dl�C~�T�K�֫"��ȫy�h�2��U���9/Q��iPݬ�?�`0uR��uJ��X�s2_�i�.����l ��ZD]ؖ�;�E<d�ozρv��f�ԉ�y|��Z՞����(�j�z2@�7���*M�1;�z,9�JX)�I0�^�%�2ow,��A�=��3[;�;`|HdH@�?��)�qW�ɧ2V��R��%��Ƃ{�Ŵ�I�a�6��ޢs��dH�2�)�#%�(�*���`��T�m"�cq�?y��We�d:a���!;�Ԧ�+ex�bB�������_�����M����M@�C�� '+�>�
*I�(V�q�\�H>*?)�"���sE�q��f��LW�t�%��/�����J�t�E�n?~� u��',Z�5�A�@�_G�pQO]ґ!z#P�>���0u��Q	�(��Ei5nlE�>L�x��	0aY��k��,��ts�����/�>T�8��ƾ 2�R�]�%6��a��K�W��%�K�7y��������[͝�β��i>vk�����w��y�=sve�1�m�������7~�����{F��e��&��[����ʩ3�c���>}�fp���0#vM�����ҶI�\�3N�8&�����,�8ˎ�?c�d��������J�������P����g�k=��ペXe+`1'/T}iCM�8O��d;	I���6��}EG"\
��4V�ty��G��Dr��7~�1�N'��,��n����*�B�����+#\P+�nd��XC��u%��n�:jE{˒6���~�N��Bmkj�:䉶)��T����Y��� �>��u8�j���ȷ=,t�	�T�b�q{��ψ/�:�$�:s4^d�<�"�>�M��G�I!t!�%���t�D���x�o�,� R8��VJ�c겲���P1!�:�)��<~�o�ȥ0(��񰁦FBa)���?)�|��.o#�jU]��w����jC)%d��G
,��I�M"�RN|��N�VN��ۥUk�e���Z�	���X�eC���*��]�u��������z��*T������DI���cЕ_T!Uj��YM��Fp]:J�"�]J�@�bcIVV2�M� (��K�0
!�SE#���e�F5�v-�.�=5m��q&	�
�-��*�������_!Z�?&����t��q�ȸb{�N�1±�
r�2<T���-��0�O+a?s5��Z-�������&8�ѥI�K#�]D�G�[d��j/���E/t��	?(ʩ�&bH�x�h%���������4&_���9)���3j��ӯ0LP~L�rɡ5?u6���1`i�`��ca�������s��`��iy�$����.C//�n��������|�����~�缤��o�/|�z�O�~��}W{�_�lr���|�����/�^po����@s������j��3'�<�7���剺] ���7�Fˊ��i㨫��tU��Q,��`*<�2N��:$�ϴ��o��y��6��a���2ywH���� Q4���%��ك�=���:L1�����l�@�8���e�I5X���˄�1T\�<�G̲1K�z�]^(^���0��W�P蜵��&���|�<���_�������E�{�`p嵧�r�z!��܈�pb�h��g8�0?��ĭ�}�v��~�jPh�����j�q糁�QVU����<�F@�2%Dq���d�Fׇ"��hzt�T*��vG�EB�X�<}��h�-"�P��`]���R�2l�L��%�E\�6���6��3�Tʹ��bLg���&NR>{�Jmb	�"?�޺΍eZ��jh�`�)���ڙ7��W^�Z;�t,��rP{/�*�6�@��ْ���q��t�L˃y�/����#�$�pcU��3X�o����H�\yI���d%n��]�L�c�*��^hm ?*�YA<&ɰg�7:���K|�Y�)J{ �!:�g�#A�h�}Cb�B��Y\���ӤS��������6u����0- ���s;ڂ�G��:���+�P�zYH���-D��=1U���I��Q�(��eV�)R����$~��qd�h�,s,;�RK~�.&
���W(�Gn�0�[<jlΰw�
9��g�M�ބ�^��+��W�Y���ɻB�$��I-��O�8�c����F�G��T�=N�d1���d���������@����WF�/�����s��2���������7���M�>Zf��7ެ�4?�=��Z������'�^p��~�w��6��7���'���r�ϴ����暅�����6�3q_�3%.,?j�:��lK0\��e	�2œ!qj^J'\��y�T^�԰,�y�i�fHx�Ki�WE���v6[,3jo���s�<۾��oo����t��t30�b)^V�-9Y�c�|N/��b@�
��WYx � �]4�ʖ�h�7���jEP�BsHC18�ݢ(���:O�^(Z9���]�������FW���~�r*%�����[:�8Yqב�?Wm�@��@2PDg� ��kPƁ���x��_��pf�������a�/8j��������u��]�|{>���+�$�]�}�Y+O��<�>���~�>rH��X�Oyy4�y�f�����NG�����^�
�����VD����z���9`A�+o*H����wth�pȗ��^��y~�<�kH9sPC5/ͨ:���v�Ֆ�*=�!���e��1�%�}���i��@���'��c�p��*@+�=���'>��J�92=)"A.��jOt�kag�i"��I�?]{�f�������5g�䣲�������v�ɋH�$�6o����wff���^u<��M� ����Y�"U����tQ"�� �%od"ʶtE�O��.�Bcp��g����N{�V�v6�'
\U��v������h�ZX^�D�f��oϯ������Ue�Kd#�+�>⁌fkk�8�ŝ����/қ���{|�|ot��j{���f�s�o�����������M.�h3}��.��z��9d�_�|�{~�T��9ÁlM ;�[�����2~3�.��9��M������ho4�nL7�e>(�� �a��OKD5-]��=��i�T_��a2��1U�h��<��c��]�:��p�m�.�6�~�d�#tC�o�c�- �RI��1�bxS��_������^�?��m^�T�J�C���Q~�$��go��4)�CG]�+p���Q��Ȁ��4���}�~D��JYl�8��!Q�3-��3*1R]ERp��*�]�	4\̬������C���&���Q��?�&����[V83�Iz�oqߦ�5��ǿ}k��?�/Fg�x�ݧ������o��]�]i>�5gF_�E�o��;����������/�s�i��7|M��ǚ���oj^�i����_�w�{������/]^[�54���7o�ݼy�]�<����0}�-���&J�0�M+�,S|\H�g�Ii��T���?� �03hos8���l��_�e��gW�E���<f��{����5�V�^$�+�#���\�����ٟ5`:��?�|<��&�xk�iԏ��`wk��]�����7~4y\ˁ�Φ�^&�>���Ŋ��u�����z{oםC<��r�1���G/�w}�]����A}���xԥ���cr5nl������o>�;�*�ɁG��$���1���:���̴�b�eBc��-Sd��x�T��ueMx���#ޙ�z[�f1I�8������_����u�.x�7Lx��ӧ�]`�5۞:u�Y[[�Ӟ�d�DĶ,�x�.�X���@m/}� �X���`!{R'�m�z s_]�Quք���l�?�}^�Ok#�&�@�H�2��Ɨ]�#^;��c��z�,���,��V|;{�,μn�h0F@-��qd��;���ge��!D_G�|��\�,1����@�����}�&y�?/;�L�� �4�' �G�0g���mޒ˧Љ�U$��r�;U֋F����8/8�S���ғO���Zh�AM/Z�����b�u$�d9�Ӣr7f0�,8��.n�� ���}>!�˷����s,���击ځ�G���-O���D�7�=���ٹ�����L����O�4K�K~�g�ǡW��F�;������=��q�n׵���f�ow=���#�4��yf�Ls�����">{��f_^\]m�<���ڙY^�K[�fڍ�����v���nܺ���ѷ�N�&Zi�hV��I���D����͊���� �O8l�W�~Z��#��J.+�kA�K�<
�Zʓ���]@ꗎ$:���pU�4���0	eK鸊@w��B��V[������ϩ�XR�s�U�\쌇H��j|���鵩�Kӂu����M#����\�*���!�y�a�!�1��9���0��?Q��g0�NH��9�x��L/�oP[���;��u>��֨��p�
鏺u��,�&�"@��9`�����<��4�Ï<�<yu�]��Tsu�V��yk�Yg/7����-}�iO��������/��/o/�n���˛_��?�K?����<ܾ���jΟkn��Ql` �U�H�4����HAׁ%��a+��3X������P�~n�'i.�B�����P�~.�B|4�ξ:��~×A��_xG��/���T���ƥ�a�k���(��q�H�G�d�L�㯳&����4�dG�����C/:�q�H(c �����c�"N�I��O��)�u�hT��tו
0�M�|�[���W�i�EQn�E�*�	�U\�*�WO��q��A�����ŗ�w�@��4�w��8�:�v����	_;=�Nhr�B@�Z� ��BJ�J�N�x�"���e�E0{��ͭ-���[��9��5&�fī8ګ�xΡ��e��-z��f���鬡�z����W�,P��9����F��9+�<���!�zZU�����U�毓�2%_}_�A��k	,�݆J�X�0�	_��b�6�o�Qf+��x}ŵǳ���X���qd#�II'��9h�`.���QD_M,,2Զ���ϔCjѣEҶ�:4���E��~���ҵ3�U3��S��W�1��xj.-Z4@˿�����$��gjp8�5M�[�xϖhet�;��o���n���N������u����kkך;.��;;������K͙3g�7lϝ>ۜ={ֻ�̼�>������^�� �������vm�����a�	ߞnoܸ��s�]�-^�w���E~{��*�oߑ=��ڒ��6$�������o�n\�-����S�E�
D"i�DRM����N�e��p��#b����a�# ��+���,Ʋ����u��Q�|��N�?|"zqB��$PɗԸ�T��8-p�\t����"��w��O��h��Η�!N˦�i^�i�cXEz���[7�Z�\7�)�.��@��#+�hcǒ��S���Mݴ�+��چ�\�QP*��ET�E���K�U�s��m�zU��Eg���N��}�[[���;���S0>sGcff���B�WD�f��o����;�Ҳ}�^����Ǜ��ls�����Px�{��|��.v������{>�D�����͛��?לY4k�����M����[�eVo�˧t��m��R�lv�H*�>����P�)�eW�1��^���2�	��ͲLO�/X���	?'�믦�t�3Ӊ�y��i��]��_�Ҽ������Q;ǅ WW͖��(���21)���X�є!؟0-2��/�c�U�1�/S�\^�O�T���z�$���s/��Q"W;�0���c�ѱƗ�C�Ϋ��d.�tbD���+9��)�k�@��t��x�ie��'�P�R^!ń���Ot*�BAc�.�uv��	Z���ie��l��n�^��5#���4��G�\������d�@���C�G�n�P�f��g<��Οd+U:�'�s�x�����
Am#‑���ꬔ��(��c�+�!כAұF���͋�i;��y���(C����J��]���`kR���/Z��>Ӿ��y��!�����/�0���i��s[��:�$E�ۗ�B'��¾js��"l3!#��X��`b��'��P-� >m�ϑ|�*s����&�M�SD.�D��9ݩ��#�"�9������;��q�3��AΦy�K^Ë�����L�e7����e���.#M����]d��}�����.�����J�M]]�@�����[>�Y:}��G��7����V�=9\,�Is���2I�/Ȗ�.0��QV�E�Efy�L4bC�A�$7	�WF«p�B�����R"<�jh��Dx
�!¨a- %@ڿ�hRJS7b�J��N�  @ IDAT8��/��MeN�	੩�tNwŭ7�_I�{�/4	T=a���0"�)�XiW���&㨁�?�6RɌYQ���S�pk��]��ȳ�z�⢄���Q9�c�Lq���.bd߀�ZPZ8x/܋S
x_w�6��?hV��3�����bA��e���t����f���²�?=��p��5~߻��<��c�K>�t�?
����|�ߵ�\�b�����;�S+����_�y��}���t�����������h�|����1�S�Xȋ�j��R[! ��?��(.�~���O��UV��t�+>.LҦ��q���8��Sy�N|�ǅ��pa�4�Hˣ����S|)X�7���L ����]j�����3��p�!&�md20M��gOUeBQ^���Z�)W����BvU�5����:x,|(�A�6�`��[E	q�%V�ӟaYE�sҗ�*� L��G�=� `�7L<��{����\�<�
Y�:�`��I��ɱ�A^k�hl�%>�.�bK0�-1DB�mc��s�n}��،t��ɉ��+c�ΜS	z-
t_�;n�$0���',���[����$�t��E��:Ov�S8
�E�)�K�[-�7X��`*R]�K�������<YRB �����u�$�B ��?A��5U�L6�\~��u,d�R����d�	-�}��e?�Z<p���(}WQ<R�`���D� ���Hp�]y�����&��;�1�O�.� ����x��P�rr�p�j���dK����ₐ�q6Z�GZ��ߢ���ϸc�k�d����S�S�� �6�X����/H�ژ�X���Z���5�O��^���H|���=vxj�y�ݫ\ �v�7��[d��)ʢ��D�[)��΅%�Ȱ*�a C�1x�g�i�5O�4�F(":�zEH	�&��Q�&
�-:'��J��r�E����hl� O1/ӥ
,o s8[�6�w�(<hO/.x�!@D,�|�\���	�P��J��FV���'b�B���n��)�yv�H@n�P���?d��q�f�[�,�8s MiIjFO�bo�V�����a��6�
����14^@������d���~�j��uވ=h��X�s˟[Ժ5'kp@a4�n��u%�~��W��y߻5�ϴ�}ə����־�s^hYO<~�}�����v_���B�x.���Q ڟx�ƽ��>��LH�����+#�qr���a�
�0��6��2�[��U��9?Y6�O��S�|aI3ɳ�1Y6�6YC��4[�l�qH�P#9A����;���_h>|�fs���>�'�c\�;��z|sgZO�>��5���ɹ��7�Ne��0�����NG,F�g�FW0/��A3?��.���8��yEɋ��m4o�H]���i�CCĺk�A�[4��`��L�H���� �ÙN�KpC�����/��4�33�F���V�<�$�vE�d���S��u�V��]�+=��t �ʥg|+Dg<TF����K+�h�[����]�vC�}�K^��gۭ��fan�S�k&�}�zpXOg�����V��C��e,��6�M���L�@�m�`�^W���L�D�7|Ȇ�M�}�稗&�d_�E�ǆ,��T�� �yy���x4�0��h���<����g��<>�O�ͬtĖ�Hm��ʹ�u΋�8����3�ښ�}\�!?�-+|�E��u����r�Yp�#�6�'˦N�w� G����ɰ�2����a�z����!Ό�K��7���xύ/���Y9QA1$�x�X��h|u-�� Ĝk�cs$kf�u�ξU��z���C/���v�'gtOm��~���~��a�޺��\�r���t����8���n��=���wp�nͷ��f{gc�9�|��l9Z]=�^�v��q�V������3��*���Cni�όx/\;�s�������?���|��7;���=47����!e�f�����J*��2�L��R��5b^g� 7[�?P�~;�މR���9�W�j�.���ӓe�PC�&L�L�ց'$Ϳ�Y���,��d��u���� ��C?:e$���Μ���C~�GJi|����(�f��o��{�H��B�PfY�����fGK�6��Զ�wY���x���Y�W�fcr�TB��<�8��:}�C���=�0�εr;y��zza�]��k֮\=����4w�s_�����bizi��Y��v�9Wc�4Գ8��u_�|�뿴�x�r�^hV��8��ޜ�{����~s�Y^=7��C�m��u��|���O���#�<�;��7���oo���.}���m�UwL�&���RӼ�	LM� \參%N]&�d>yL�I�p��t��yN��e���'�d,�!KW��Õс��C[�jڛ���=�n�N����+3-/�4�O��:;Ja�&`2�c��J8q�F`��h�&H��"��O3���{CQރ�h�HX�(�;��%[<�=Z�*/yQd�C� :{�^Z~���"�n� fߗ��IB�/��d�ðL�^D�L��K�F`�H:]�Sx*$}����3��K�X�/^cM^�waG>c�<56bP�E�����T��hZ̸\oMU�5�nm���tkB2��&x?�����o2��2ѝfc{C��+��k{I��x~~:�Xp�Ʊ������X���λH��&��)�~P����D�io� M�\�p�Za���{Xh�s���s=� q�h���S�"`~i����v{ͳ��G-���g��Gp�WB
��]����1��b�3`���BGc�� <�L���v{gSO��g-|����i"�F���Y��m������Up��E�CN�0%��؃77`̩zU�~�����B��F>������ ��b�Ş4>�$�_�0a����z�Q]�л�u�CA�SO����g�+�;li.,/�>�[�9L'y�����ں���ikk{t�����.���"̃�0��%�pVn�Y��@w��+v�^�}~L���9�!�e�g�?�<���������R��������������}�zz���{rڜ�]�$d�ńk���g����al/��,_��`�8`c�`�`�H\2�E"H(��Z�j��N�==�3��ߩ��?�]d���>��w�+�:��N�:u�W�����<��
�F�!i��.Ҕ����a+l�	~�e�~j����O@Zx�=�Ǉ�!a��s�����@�,|��Ć�?	H�
K�p�n���	D��0C&�D���"����ڸ���
M���3�SyŞ�8�r�	>I�4!��[Y�����h�	1�J�	1��"'jÛ�Ϫ5Y��^�����A�Y�0�2Oӓ�Cgf�tV~�uE���S���l(2��O˯���(V�\ԩA�V�Ȓo�^m�>�|���k�����|���˝km(#*M��DݠkZ�^y�d����������ֿ|���g�r�y�w�/~�&?XNܯ���n�+��=%� :�i����W��|�_��(�ށmn��fh,@,+1§n��W��#�
5J�Y��\�"?�+u��kwG��q��
�~���1N{z��/oF���Mî���[.�$4���Hw�t
U��1sq�Ҥ�U�M��@�~�]4�Ss�,X'K���D�`�.X��ú6�IxR)4�L�Y��K���1X�f� M�
�,'�Gp��[���V�"�p�~���s6�^��,�P��nc�8��c�2˺�v{���y-R�-,����g��Ѵ�Z�7�����Q�Ư�:�9&��"*X`
:#�\���Hi��6M��
`w �+ ˨vm�am`u�0)������arx$�:Ȧ�wp���{	��sp�8$Z�z�,�Z��ؕ �t�N\աy��X�[����̩���'�� �7���������A�ȩAK��ro��ާD����/�W�����O�
tc���88������g�£?�3��eT�2�O��d��P�8yS�>�Y�F=Jh^�`�0�/��~��hzOIeS���iV�tտ�� ��+1�K��&���y�z����Y���&<h� ��ȡ#h�R��Ϭm��]��7�P;���O�l0'(�"��vk��˸Q�A����fMD#z��F�e�����Z���d�-�Y�����F*��4̸XY���m�~�6,��q�OL�d�:@)K�H���MD 	��x*��V_�|�F���C+Ӎ�w�S3�9� eͲ^v��i'����v]��r�)��֪�K ��_��J_��>5Ж�o��?^fh*�����mMˠhUpE�x)3�c�R|����W�b:%�ȉn�hf��o���U\>� ��Ϲ����QJ��`3��U4�Cb2���'K_��O}Hf�֏PF��X��}�c�<k~�<�8�����;Ҟ]^t�k\(pe����,[̝��a��Z�*�Ձ,�/��P�w�S�1O-x!����g���fճ�4��U�<��{��g��
�Ѭ9j�z��\��XO"���kt��9���Q�{���?��й�T��;x����sT.�{���;m-����?�q�K�}�۷w�=�I{���t����I��.6�?����*�'_�7o��ب���а����*��~)x�	.��8y3�D��q"��n��K���j�+w��1纡�E�v%gB~E�tu%sk�~�2B�rTMW}.iΜ�kz7�;�I�@aa�c��R­,jL2�i�U\���.��O+A�2�Z�����(�|�Oh �>��B	�V͂&쾱|fKݶަ���(�����q�j�Ѡ�Kqb�9�F�O�ah��[��r�b'8�i]бY�EP�H����]�9��
�����B�H���܊�js�LQ;�N�����HHI�6�!�}hT���Y�,�;+�mIڪ%-�*��Cܰ�&��]���E)�$�ObA��m�xt�P(s�o?L	�Toh��]4����E`e��%m�hR "��@�Q�V&�/�8b:��W���͍�z��Q�����������L1��ּ�W�0�]J}��?)�W��>A�{��텴�n}�W<�W���e�+��&�]���-Vvs[��U�fiY ?��������G*_�G����E�)\�!��L��Z�ÍI�"vPcaU֍Zq�D�Ӽ�^H�TFK_U-/�f���r�SXz�xr��
�0�ˤc�.�Q(�]?���]2���CuC�'�A��
�����|��;�ı�"�K��S}'��$S,����j�]�zZ�%VO>����昙��� 
!�y7|*�:!f��ɦF�T�e�@h;Ʈ~��E�V����u��^���d#�)�"G����"�	�PVn-�m��2���G������~L��j����2��Ԗ�Q�>����Z�pZET��XhK�'�1O8 ��iq7U4`'\	%��Y�ꂝɦ�ip�|���
y�<{"),,�.�y��d�R�"V��9�-VPRF��
���5@y�X�4!͠�+���TW&)M>�t+t���B�����F�a-s�Y�y���)CgWUj��ZZ�a�U���1.9[��m�R�(D5�6���Z�MCW�7Q���J����������ʿY��IR�4t?X��*qu;(�0kg2M{	�?�i����+�H�wt�ʮ���F.�o�'�O:
˰����.�������>�5zF����F��ϗ�-�|��������7��z�~��W��	���r�_���/�L�7�������u��?�"w����/�'(?�c,'d�d�`h3IB_k���qSzE��wf�.쓝O�)�˻��1No��`���1,��/���y<���a1�|�:#r�k4Rw�Z�ѦXtF*])bI���MO������n?�ٍ�?y�+����0FI����l*s�(��ZR������,�?-h`s�y����݌Q,�ё���V3��g�'�{Dh�L:c�!Lִ�T'�73,e�r�<3���R��ܸ�Md�z&��[\fGK����-��k��?���7A�����F��g$~����I@@�E���?�]*��/ju`nB5i�K���є�s�����$���<V[F,,睥�+�� (W.���,j��&H���L�O\��l��*�b%nH�e�G�v��A��gK^�� �6ɍ��e&�Sv ��bD�┠�nk{�7�Y� &�ˉ�f�G��1=�rG)LVִ�;�Yֲ2��*-Kq���~B�WI�'x����A��b�5�Pե���R ��l�Y+�d!�,��Pk��Տ� Ȓ�i���̝��}�-8�j3���O�-�V�0��S[�lM�0�5VhqTX�!`���8��X��/�?,geF��$�M](ܫp�%�'9�.�,����4�^/�DC�f�d���K�8��g��ͯ�aS�� z$Ѷ������\����܅�g��� rw��Y�w��0�N�XrT�ث$��+��c%'ڤP`�m�P=q�r/Ga����$���4�z��ʆ�K��e� �n�uq����X�%�����]�xl�"
ȿq��μ��VW '��m#����e��E!�6 h��q"��_D7l�����Eڪ�u)>Y���3�;�j^�6�%7��-U��Su/�p��q?�I:�Yu7�2�&�"t�fzqÏ������|�?;Qs���rC���>r�k��]��nT��2�����o�����	O�'Ϻ��������v�$����Ĝ�.�QwQ&/��1�ݕ��%J�p�#G���M��aF��"l4/G�W4#�v����ǋ��,6D��ѭ�������$A���aAW���ra��Xw����_u%W��Λ܍�/���e�Z%�>��nN�TV��舦Up����|�aj�����`V`.Np1���|F��������0Af��J���F(��'�c&�������3���V��Cz"|TR�PqilK_���H�((�,Nt������ã�zY����#��l��gY
͠����ea�D���R���4.`!�~͖�g>�6A*j�`	1�@;\-�<M/����J'�Z!�3��L!���ֳ����?-��L	Y[aV�փ��^����[����d��|�	Ij�p�9�N��_T��z2�ށ�0�S��ڶ>PR!0�q��Z�6��y˗��Ky�H9�G�#�!/Joq�4g,�<���\yH�ͪ ���5�J��. ��~�K5��3B
�@�X�'�Rª����1�n�jyDǒ	����E����Oڭ��31�������J�� R�S���`���xU}��Q
�4�v��\k6�N:�AgT$��x\X��G��K��|L�g��F0y[�X�������z���z��Q���f�.�H r��z����prT�q��s�B"r)�!R�YL�.z�PsQM����9|�����\^���(��ȏ��+�|ٳ.tQ�,��2^]�Xk��1S�=]́ҡ�Γ	u�H���5���Y��M��ݹm<Y���+��Z>?����R86�c�X\����&cOչL�Px��@����>��;���@ȓ�1����J�CdG�r�w��SYJu��)Q�o��Kic�}�Z 	�:=]|C�35�Qc�vr��6��@��
O~���wN$Ş~����=���)����^���������������z�{�{�����w��G�t�b�TF���������T��s5����Q�l�)yu>��c��f�O�|"��`���Hr���ad�֍0��o1.��(X8"Xė����/I��TD���ّ�������B�n}�j`>��k�������^pWr㽧mw	���l�~@���U�B�g� eI��>�e1����˒~��������2?K�ʥ&�ɶ�����⌆��JF�P<Y��g��+���0��1�/�e���r�*S�4"��*F�*'B���yf�f�_���?��C���&�җ��E����	�I|y��'���
��F�����"�˨F���(Κ>M�|x�~�3�o�f	��t��O��%�l��wK���f�k��@s� S��4��)h��_���Sx�e���#�\@'3+CY8.8����7���0KGyj�QV���� .���j���AnIC���~�L�`���(hO��N䯴�~�,i�
B�	�P����=_6C����X�)aq7V/
Q~��*�ŇG�t�H1����I�_�Fu�̛��:!�`W	Ð0*+��Hg�,�A>�rX�1bI�Onl�M�R��kg869ġ��9"�� ��%�T�TM�#!}����c.�<ѿ�m�:Gޫ(.�^�NN$�s�ҹI�fX��:?\�PYGN�� �ҰBX W�|�f�
}�Y[s}��d�kӯr�p��y�X�h₄��y�t�Ã��A��&�q�K����
~Afq�l��0A��֨�*ԃ� ��C2C�CQSԇ5&�j�3�
\���Y��n�!4�7�653i3g����t���x��D�y�d��y��/�����P<�˱=/f��ڴ+�ر2��f�g#F�W�SxuC���@��DH�g�h��7j[u��Ҙ⟵�:/�)R��*�3d��V�2� F*���~DB�=���C�ݱ�|�>�����-U�׍�&y`���7�9�A{}��N73}���_�וF���νn��j,��j߀�7��8~��dhh�*~��*W�_(K�U�,���ղ�r�^��?��pi8����i�~"��R<fʮ�N������;�Xl2!Xe(J��A�g�gg�Ȏ=�4C��c�P~��^|��O�iY���9-o����§J63+upI�� �?���Ѳ�jUY+F
`�hj��ŷ��Mȥq�3Fv�c&,���&�� p���^b�l�fy��m�`�`�~1��*��L��=���*� mU�� 0iy.�cYc��i�ƴEQ��=|/[*|1\�BX��zxY�"$�<XZZX	��W�8c��ʥ*���4w$����	���Q^ �S���r)Ĕ~��޺��CH��(����W��Y}F��5�yP�R�ֻ�����1��/DYV�K����J��o����b�?�����RJ�Vw�,��q�Or��"i�g~:T>���S�յ��B^��tc!<�F2�#1+[�B��GC�&R�W�-��Z<�l�:��jo�0C��Rkʪ�M��F'���Ǣ)?+�<dQYU���J���t����Ԡ��0�+��A��% 7v���h�4���&7Z#�H�b�� ���\�g>`��M���',����
GH�Ŕh����� �Ԙ�t���kx������Y�7�һ���$ĘG5F�V}@t'y�b���A��ȝ�9pj��pT�ct�-����]��VW�jΛy���8����\	'�����z�,R�2�5�Հ�J�<���\ot̹�Rw��	�l��e����Bm�SjP�thc���M��i7�óK\.a[��<����Z���֕TwVݒ_���y��L�Ɗ;y�]n�����B�Fǁ�Э.Os�
Q	�����j���ȁģ�ݣ1��N/���~(2(t�0����m#�Ԓ��l��t��COb�U����hs�[Xpã�8�]r�t��ω,�|��i���{���f�	Ί�\appn�B,�.r��@���d��z�G\7���*�Ij���d�_Bf(��?�$�Ų���ʦS��~�$\9;�/��=��+\�1��O������oM�X��y@��w�8"�\�=α}/ו���-7��	�;ؽ�E�J(�8鑃jK��आi}�>���k ��* g�/�Y�#�E��w[��#��oK8=TC/&ZEn͵1F0��ą@�!}�g����rPN�t�;L�6�8�&@0�N=/�/�����$����Z��cVi�,ۖ߈?W�<�'�V��pN̓=�krI?`h�'J;9R���Y�梶�\���WVo�-�Ԯ��"�H�,?OY�X|����9b`�k�֏4�/�˺�p�2(�V6��pg�BJ\AY��L�d��W�[�+�~���GCu���p��<��ư��.��n!��P}��
x�n���reR���E�0�O���b�K�c���g�knmH9��#�f�L�Q.��Nd��(�"���F�,�b��!Ǣ��T��f�P�\��D�j�*3f腖��bʛ`�bYl5u���"k�S*��6	�+�*�UJrpH�\�L�+�Z�#)>�
�3G�c[�Z_9�gk�&t�eG����@��>A�x\!�l͔�Gu��~-�,����$߉�5��*"�E��@�LO��gNB���*u$(�p���m�I�N���m0 �;���������ғa<��mٕ��@�>�J��}v�B�:���.t#/$��Zפ��m*7��Ρ�F��dmr5�s����fRF?Vcq��v�r�G�yʣ��]x�a�>5�T;���J+�W���'��q�,�#����(~�ᘒGߩL#є.I�=id��!����T�ĽT�@'�~:_�*�����R=�Vl�>E�Wj��%;Ԕ���U��I���eF^��l�.����H}j�;�*y,@�ltP�A
���"Ԓ׳W��B"�h$K��Q���¦��]��-��/�被��)2S�sv��_ތ�y?���r�O8���
6��x�f�&{�_���ad/����x���fhJ�����0M����N�.C�� ����X��NZT���U��
�b1i�|��'�
T���y���gpJ�<Lt�Ov}���5�|���r�F�M_>Rj��(_*�ʎ����òi85�4���J'�� 
�M�g;	�X�*5d�3��eH�jA��ur�[�W;�}B���o�-�𐅐��� g�P�C�-w����������o�7Sap��a�t|�GY�M-!�heL���l^�a�,n���_�i� X�� ��CV_��(O�6)���	���je�,��_`��8x)����:
��7�g�� /Z��X3)�D's1Y�,ߖ/2(��71����R�Α�mz�[��̆`�),�Cy�^o=Ey֟�b�+�}ʋ"�e���R���>D��#8m^sL����݆ ��bi>SrjK_��>���)�Gz�tz�\�Fc1*
�٨��GOR���i2|Ѐ�����^ !ԡ%'B$Գ���Q��*��%�1�1�	=��j�N�ԏ�fnOG��Σ�W
����c�S��U��n�������`5�z	���Mmq�w�W�*�7���M��.8L���Q��匆���#��"7�!a�"m���Hzy���@�f�<ˍ��������cȍ�������۳m���̻�����²�a���W Ҥ�b���R���q��f�/O�̖B"��C�C�mk)�a��S�9�J���ϝw�%.D�!�5��<�9Pu=��ު-#��{h���1��ЗV���)C[�\<������a ��qi�G�i�(B[��g�:�x.H��l'hTQ}pg�!���pC",F��z���f]Y��t������4�0!�3ܹٯ��[Mʬ���؀#6;�LW7�f�ms߹Z��]}�Wv!h�\�2���̕�]\�*%un�qŊf"�[
(U�x�)���9R�Qshڟ	�m��T�B�>�ؖ둶n��g���p�0�G����*,q���9�HԹ��3��&�^���h�NK��`�H]Q4�ԫص�#��r�J�D�?�qCui��j���ab���EL�������r��)|�Q�l������R�14�ff��kD�l��F<-mr�Y�����tOf}�e�4�:uj��/�{���D6*cr�*O@F�jO}��B���.�� >�̒5�ܚZd��i�ɝ~���=S��,,��5�l��iʱ���|�!ۊ2�rǈ�F�˕#W�����&�`�#Sڵ��H�2I�V�<a�(
Q�k�X�G���\�'�4�yf?��r��ʯ�=���EP�y=�+�"�����i�i}��O��t����_>,B��?���!0���l�|�^�-Ė;�1@Z��c�ӒyEw�Ov�:^�%o.6��n0-ߝc�3X�r���!!Ci+	�����~�����K��:R~�� b���%s�N,z��!�Xv���bFa�82щ�O�WWP�wí.9n~��C1��qz�2@1�ց70;]o�?��E&���4-"υdfv���Vs7�A��k3�j�r$'ޘ.�K�U�nH&�$]ć�C*���Y7{�Qı��4wIh��æ�gM���w��ew���	H~F�a03���ts��P�Ha}5ل�ٳ{��V�1ZD�ⲛ�I2s�M��('�r�5������w�ܭ^���O���u#U��� ������dqy��^8�{z.�'Ξ�K:鮢T��J�ճ�:4�{�unJ�k��ah]$��U6���m�ꖎ�q�NV81�[|R�)�J����Y�U{�%ƜTC_�mD��W$�n�C\;�uʿ�b��K�g�\1/�@ w���olp6ь��՜�u���ptIF�P7�u�[%�>3M����;��5�i�N��q>�'�_5�E7��� $f�Z��ߖ/�˓r�4�¶D�!�|���ᒃ���y)�_�~�D�C�H[�4�rDmUƢhWF�^�X�Z���k����b�,k7fq�%�I��ͦ>f}C.[Q5-�'�!�Y����V�pVyT�j~+���o}[����o��j�.��oTW�:��Q�@"�/�CpR
7u,E��J� Y�%q�5���gZ��QT����d?͢��Oju��e�S�(�)cLL���M����[�I��=�/F���AZ緬�/`C��L2�����l���Y%e�r Z�b��a��$���5����X��e�#�Ӣ�hF�`��|�j�!/�����4V�W���/� Zp6��6ֻ���h7�K$�T� �YN�/C]JW��TtU��u����n��g�(L�;g}@�#��0��2�4���@}��L%��,}ć|)j�	���%n3	>-D�d�L|�V�Ұ��N������Og"�C�d�6���Z�0�Ve�S%�L܍p�G�UW�٠@Y躶n�b�et��bބ����uY��#�D�;����nر�⫊��ج�*2<�,Լ�ŻbR�='��v�Z�!��T��ʼ.���٥�x�� c�5u��CL設��#(�'z�*v\8?��:�pҁN i$�O� xB��r�;y�Aښ[�Fܦ��n�>o��;��G肰(KP�TJV&���r.��'7������>���v��,͹#cnej֝��AĎзD>W��0�)?�B����!�2�z����_u/~��ܫ^y�ix�N����׏��*�.p<��H��SU驒ޒ۵c������KKn`|���U�;Q<�3D^I7�,l~C*n�GH�u�u����N���&�.����z:���yZ(��L��\�kK���{p��q737O�x<�����5:���SqSr����(�������Hap�C8�CT��O7P? �����[z<,ӏ^�����d��	׃�|0QB>��s:m���vW���_x�k�����o{�+T����q�"��%�xɋ ���LZ�+@n�_�k�~�+];��4>���B>ܛM����F#���t|�q`s�1<z���o�IJ���eW�`Rr��������˼/�h���Ʀ�Pӯ��5� [��;	�J�� ���fS��+ѹ�%�Vm�8TY��X�
�����\���f{����rx#�{98�+,·�Y8,��Ul��N���f��Ai�N��Z�B<�����p*|����+�iG�*{H ?ß�/u1?ښ~�S,����=���53��|xL�L�/�~Z�98���oI?�����y9�ϣ�)<�?Ƌ������2f�m� }Y@p��!N���N7
�j��L��)�?�3r�?� ��9��.6�>e!'?�/_��h9##1NTĥ��,(���z!n�G8��f�;��	�Ȳ�VЎU�.���&
6E�16��!x���?�B���x� /�7����q�]|as���g�+-���k�_���\75���͹�������Μ4��Ơ��A7wz��x����	�Eoz�;���|�7��H�{��s�����#��>���^�ܧ��q�~��tӧ�����w�M0�X���YOI��8�冟[��
�U����-��;w'�(���x�m.��:�;~��qd��P�ĭ�_�u�d��uOx�[�xl��Yw`�I�W�/<t�#���[;.�-:�1�F�B�!:eXW�f�&�ȭ�Vѫ��'\��[f%B��>��0� >Ո</D:���:ܘ��[[�� X�sS�y2��8zzP	�6�䈒mU%!���bIjk�����4+:r���ԍ�P��Y�@� ̜=���Q��^�?5���ħ\�8N����tX���O�j6ys.<uj�G�#���P�I&غQ>:3+.�!F�:�d�E�+���+�6.�U�:B?t�^�"�b�<qE�s���3�R�+z�-�<ǿ����ˮ���~����_��k�0�߂��g�����.�F��mC����
6HGC�s�(=]4���1�4ؠ�ۅ��?�&�|����/'oW��4��
+�zy�s�qD���g�۞׸�.��NL�+ĴrKG���zer6L|t'UA������P՚PV��/��~
���ǰ����E?%�BH�~��Op�?�g�����dv��UM-�e`�ť>��p1� �S�m�/&����F�#����5�N˃X�+�����ʏ��IZ��X�)�ܴ*�BÇ-���|!�����Rx#TL+����I��8!nK6%�Z\�MZկ�A��D?槁�ڣ���J/��>G_nÑ�3��᨝���Bc�O�o�^�'�?->yN� �8Z�b�c�2b���N S�,�q�V�օ�h�v�S?|F�*SX|��~������
m���0���K��J�����8����pA[�Xt�[� �����Ӂ��˚jb0��ȇ�gı�Fn��z ]�k���@���aD?�M/�4���V��6?oڤ��%�xϱ%:|�\��qL���溸A^���9�lD�f-X���<�\��:����ݱ�guj��r0�$�f��H֖.��s������)��u?��������A��L^����lδjS~��7���Yw�ܙ�S2���5����m�l�9r]�X��5^a�#wCo8u�hr�������u���!���0���}(�����'\�x�����Iwd�~��\�'�9&פ
!��L�^��Z�<I����FarnQB�twn$c#{���HCC���|��d��\@j#hntt�qW�_��kImB���s{��9��s��Y�#d="�}l\2fI���_��B��ۻZ��ᢪ{��9r�=ļıfO��ב��*U�M�OCjQ�suݵGhF�E�d���By�v���k�>�-5��w�����s/rN��6%�nl�54�s�Ho�������$p�c3BgWOr�����w������k����㦣�.�ܝ��[��M��$�'uw��߀;�<cf��˟��u���O>y�_��g�OY!�`<�}���U�u���$�?FS�.@21L ���%�cN�)G�t��P��k�aL��B�9���-��=���c8a:��	:�5�V�K}y�ў����p��ь��t���<W�P�n�W��[���C���u�9��ql��8}a���#0��fpmu�2�n^
6�E�o�bx4cx�a�M��X���Fh�Q��v�S�ZC��w
m�	�}�e�$�Z����"��?�������볎aR3͆婕n�}`,\q�]V�P�-�2<[|[e��ь`y�e�O�3�X�h��M��O��V�7�K�+�+ڿ8}�}y<���3�G3����ݼl�S�ɞǓ��N����p�xK��qD۸f�=�Vi�>o�^Ջu$�@t�ց�	5�ޜp�3���	f�&�Y�N�)�  @ IDATA�� $@ۿ\"n��%̗��0�\�m1I�����"��9�0���I�?;?!J7� 1���!G�PR�.��ū|� ���M�xfΟwu���%��;ȡ&�pR"h��+�:R�����`O�,MOZs)?��
k�4F�c4�N~�E{i��w��A�(�nfi.����z��������{���&{�V��~�8d��o��z����u��K��n��	7w��A�Y��(�L������wp�鶕K0��F�g��t�~����p��ٜ;��g�'������D���z�y�vÝ9�P��ח�8��N*��1V8E6�I�Zg��o�Ź������M�%;�mC�sG�p�{�k��jhF�::�
����vK�:����g~�� n��y�mwW^q@�n�m۴t7����:��l<�L��b|	av�6��Z����������>������~�{�>t--p�	�#e�̓��^�!_��p��˿"R�o�6lTC7J=5���҂��'����[�x�Op=DV������I�r#��o��8h$Ĉx�*��@E�2@h��F���/�ã%��~Í��߸���ַ�>ݺ�}�u��u�s_���[ޱ;��W��G����y=����<S�O�}������?{n��m���}��sU����U�P&I���"�l6���+u���raPj��U��Û�χ_.�\.�_�~q���mA�{7l�u��,�
� I�H6`�V���h�Pٲ)�#�J���Bd��X[���c��6�-3�o7-�Ŵ����=q���=�13]Lm?* �"���^2=D���j%Дxk1`a!�
Gǲy\���я&~݄aP;��}-�_���ai1���(�h�e���ا@,�)x�;���]�4Zjn�L��7� Oni�s�R�qf9�����X߸C���ha���0�TuQ� ��S@�	5��"�m�D0KW�1�[� "G���\Q!j�G|-�O�A�rC!���]�(����O����G����_�m�'��?b��T*�?3�`��S}�t(ibTR���:U/E����!!����$M�k\SE jO뾖.?�S����Q%��|g0��1� �+@듡�2���ѦT�cqA@��j��E +&h���7s ���Hc��3���A#��c�bW2Ĥ8=q��M�ӎ���,�,r�w����\�G#D��@@�� ���_�x��s����'r�i���l�lٗ��ӥ�z�ϟ�4ܐ����^��{c�+J��}�%/�qw��)�����%/{�C?�Οo~������칋�λ�
��6�<��O�_��W�+������%P����6�g:|��<(�f�j\��aء�+��>����?��~�WW�e4@����I�{�!��p&Nsd��)�ep��[Z-!>��d��+AӶ�XF�eM�o�w�j��'�=*�Q�OU���t�=�����K��h����3����P�G��1�у�톆���S'ݧ>�)d�jF�TQ_��!�d�$�{c���Ӟ�������h]W����W�������Q�Yr_��.w�o��|���,&���z뭷&��F��_|=��m����p�c�e��7�,���q����`��%���:ʣ̃#�]��0�#��[��P�k�?�����^J"q�ü�t������t�sSɪ�#�F]u�[^Zv=�W����O���F��~��n�w���o�
(Kn��������9�{wI�%�1�^��s�8�?8G�d�=����Է�J�W�4��݀�iwG��g��m�'�+�f�!٣>N��aѝ7����G�V�9g*�����:4��~}=nxd�M? [�F��
��v�������v��7�fƸʩ�?kL}�?��7�`�~���S�O+qZ �P�ї/�	��4c�>����r������������o���,����Ȩi��Z~ඦ���a�+�����75}������fC2Tm���M0]�q+}�O��iu��<o����������,������9ұs��pY��KS��c�+,L�!9�-��`Q@�n��_�/X�M�}c�
`5U�T^�^�?A���D�������m��$�b���װ��:҄y��M��+/�@�r��^u ��<'��*��0�j�Y��p":��\�@�!����	�B ���f���z�����]����<�����+����^��L���߄�l����VY4Kd�"?��Os?�3��}C72��3�n߿1������z�3ݾ]�n�gA�����A�i���oys�9���/}IR[����_���\�����܁]���8����ۆ�Q���!x���:7>2����7�[n����w�!�B�#��(��n����<����je��&!�#$�&[}���̦�n˺%t�1DC��޵�u����h�M�]���~�M�r�۽��7��j����>h�ǵ���W9~���{ݓ��d���Ƚ����b���&kVA2S��95;Wn�>|8ٱ}�q�N�8�l߾��~�S�N���_�~��?��~�����o{�;�>�I��:���������Z��M�Fm l�Y@�Gn�v3i&	�n4�q��:����~qzJ}�A�Q���ܜ��"G��a�D�]w���(>��&޲�Gx���ήAOM?��J���<�QZsCc��¹��oo�K��'?��w�@A��6x����S�+_��7K��"�:��5�6l�1��i˛?�Q��� ���[+�j�IǶ`������ϻ�[���R���[}y\�����C=}��	o"h��@�i(�0��&-�<�lD7Ъ
�4,[}1�Xc�19�$	$�O��R�`��^A��� 1l5c�,�4�[��,}��,W���.���v�'6���1[˪	�m �4�ڬb<�5�hu
��K����~����#��u0K�hf����n��?K���t|&���/M�
�B`��F3K?��Õ�G�Ң��4{
����.����OݏH?�����v ;Q���h�`�~�IW$��*��\����\k
���oik�V�C>b�{�W��~"��?K���o;sG�1i|�O_�nnM,�Y�S[Ch���=�a�K˞� �?Ri}@�X��l���l6�@jҟP�B��S��vs�v^!LS���FHKU���/�í~)�)t���>�rg�ȎQ��ƯLoc�dķ	�}JN_Zɪ�E���OG6��UN)/���<ܞ��sI/��E��pFe��,�)q.U��W��?6z��~��@�{������:��o�#�4�"6	7qa#Ѵz��Yw�='���4�{ٸ�t�y�c��>�1��6�Ru�u��%�~����Ԝ�č�n��Fƨ�j"�
�k��ν����+~¿����^�S?�-�!����87�x]~a���ь)�N�V�/p���>� �+e��s���2%8*�#�����t�X��0�+�Z���&�[b; ��QZ���p��*�P�����(|�!,�{"��Α�?.��=:��K�P IC�;39�&f�܎=�F��Z���?M�sn.��3U�C���;v�I^9�vcCۛ�!78��P��=�����v��q5�2O�����|_�79u�a7�N�~8F���1�>�1s�^�j��w��߶���}��*Q�%G�&\uǶdd�^7r�`s��7xhs��a����
���׳}�-#�VCX_�����:a�O�>�:�i+w'�Bn�k<)ѯu�Mk�F�;N�2���bLN{���
��s��:�S=�Q���¦�s�;Pf4�����]X��-=8j�Z���/�����P�E�Kژ��h~��t`c^�Ƹ���1�����&�(�9�EP$} �/�l����.�4^:��<�£;�k�;��F�h��e�p��2�b�7x�P�ҰMJ�_�>��SA<�覦�����O��	�;/"�dȹ��`s���7�3�c�bn}�?o�ygVŋ0y{�aaFk�#�G��~��b��nfiH����!�nu�5SH厦�
L�|�y{��xF�cQ<�E�h��2#�4�Q��B�d�gN~���K�4�]8���b��� R�%�',�o���,}�=��@���$�S~��c���J�e�6�Z��q�~�b��|[����m�J_��'�ǈ"��c��	[��ى�&����
"��Zv�D�P�t�-�,}9���@� �	��M��4MZ�0� P�gi�'�Y�щ[<r*I�\|�I:�є���8M6I8[�� �ַm;�O���#�ldl�@:����:�D�_��;S��>ZwA�<ͳ !1K�"�S���b8G`ia޿�G�w���̱����7͕z���&��e��7y �;��&y����߹g���ם�������t���㮾�@gݻ��
�ׯ�nT��@���o�i��t=p�i���D>�[�r���'��8p��q���l���rT�kfn]=,ܜ1��T�`]�5X]K�+I�������vZF
b�o���l�
�*V��P�LȰ�z�kV�"Gm��}�T������.LO�Qg��Xs����A�5G��q��s{}39r����c��_�B��%ݒ#�K�0����}}��{�����\��5��:G�g>��(�5�	����F�� ��C fM�����O���������|��ǃ�~z��"���T��P��C� gP������1Pn��q�����:���I��pſC�J�4��U��]��a�0 ���m�)�U�U��ƣG4����ɺɺQ��tΝ��F�;|?��s�.V�l�R�.�`G>��ǹ^4�/�W����Δ����DF��7O[B������U�4�D�r̆�ԝB9?mr�NG�r�Oc@v±$��a>�����"��L�),�7����_��!�MH�U�O�-hOCr�du�&7�BZ�]���J%!tG���&�[(��k���!��v㰢i���Ga�	
+��C� �E�R� C�ʜ�Ds �0�X���v��~�W_+���?_6C 9KW[���ڒ~ In��F!&�2�X�IT�t��Ǹa�������$a ����e�`PÂf@�n�U��'J׃Â��R��G�pfȦ.[OԘ
ծ�>-@��x2�B���&��*z��C{����ǜ��`��Gi�⭐O1R|i��\:Gт�%X%�%�b�����0[�4#1�X��g�~���4&Bk�Ck��RmkQM!��ťlۓ�y���x��%!�bg��z�1�H��[C{n�Ir}�[3��O��`nn������P��7�x\dA�,� 4<��:� <Kdp����)�5y��_���X�C�VѬ:ȏ̴X�z
�� �/��"EȨ��Z_4)c�n����11;�t��Yi(��f!��Edz(Ox���f]J��΅2*��kWu e��0|}}G��m�q$Q�@�5����ν��IW�p�q3�
*�,��G.]C#�k���@(tQ�.�P�Y����5��or���n���������HA��Ң{���z�����[��vo2:�$-���>s���n��?����[<��D�x�{��3Ia`�'�xm���r_����m_�����ݓ8B���i7r+�Ο��p$�>���ѣ����B�'%��p/�LG�������pY!�:@Qcm�͜9��k�;���E��m�Y�%�k�������1�����\��;�Q�ق��E�����]���+����OX�!���P[�������_�"����Ο9߼��
v'�+������m��a��"*��+p�������0�۶m�����iA��I;�(����s�Ւ_�y��x�M�o��M~ׁ]��:�md����9�Qܸwt����ov�t'c��F��2��2���Qj��lg�Ϻ���x�+ wu�<��c.�=n���Ϟ�lԍpZ�^����-��F�g�F�/i�A8l t;���(����!D݆9�[\���Ƿ5��Got��7�
�'h� �����?�z�����[�����%����	��6R��xg.���%�U����.P��I�j�~"�Vmx�G6X/A�?7?bm��)�G5�F"���;����Eْ �:t�g�5i�Z����(q��@��-��r~�Tf� �
�>M|ў�`\��;��h��ߥ`�q4�_
&�ʛ�p����_H_š<auyd�ZH�X駎B-��F��d�̒�O���D<�h"���Or9��b�������_Ւէտ�o�iWŅ[D�ա^h��5��~cP�k+\@��N��g�҂	�-���0q�!��/�����3B-d��R0�d�2	"���	_�tir,4�������.n>qa33�(���Ǧ�S*l�܅�ik.�Ѽ�L��d�9��^!fW��D-�,�'���'#�����Vyȿ�?,��E+	�t������*\!Y�М�v����@���FQ*�SW\//�x��еln-��5�s�v�k,�DN��[Ԣ��I:�^��֥�ϯ�.���F��۩�&���1Z���2DA�_�F��fw"9f)��l�Z��d��.��iu�W��ϱ@��r�}�'�����C{�&�1=ksn��Y��_�E�������y��U���b�*��Wr������~�M����C�!2E����C��L�&�?���0ϻ��qh\�@ K����2���xЃ��/J�/Iy W���,�g��<U�%�s�w^�Ξ�/L�;�BX�]�((�s�]��Djo�
Gl�#�*ς�ADl�
��C,��B�RW�(�%s3S~c����,�+?�r�����7}����薸�v���\H8�������׿����O|z���O*#�2h�N�U��߹sgB;�d���G�]��;w�v;v�I��|���/��?ppW�E���ɽ�r#��Bx�^�b=p�x���{����C�Q�0�V&�F�w�02B�%�F�9�͝�Ȑ+��(D�&��2oؕ�EX�y	��@�^����**6u�R}�7c�]ی�'Jl`3��*p��=Ȼ�3�r��~&q�>z�
����� h�1���]p�x�Ӓ}��W��U�7���<��c���W�8n�-j"�$m��Zѳ�FA�߁-�����Hi��}�8��c�kF+d�|��D��#S_�O͌@ʇ`�O���M_�%	D��ÚB"�a��N���	b�L��I�dզ���.���V$����=���yw��a�3����g�?�cXĝwG���T��+�֓9��2a����3���b�m�8�L�0]�7�����d�մy���b�g)�@B�Q�rG��ix��o��-qŕE)�/~�ng�Č��0l#�l[Ɛ���qv��M�3bC��MlbZ[(D�sLf�ʜFF�%�D���K�i%��\+:q�1�p�3sk�c��(-1�"�$��JF2)�B�%�ŵ���A��w"��ӄPج�~VvMn����b	�����D�/�$d(��$��:#��U4xh(K�~m¸V/6?s���_^XZ��Gс�m�]�u(	�]�wFS�̒���؅O������{wq|i�E��������ow���D
�8%�	Q$*3 ��@�n�5)�U�M���'hֆ��LNG����˗p6{v�u�.d�v���e�#�8^C�
�iQ^�6d���Ԍ/@@�+���j�hq�-o~�����?|��������nu>��_�ixr�8�A�-.%�N�ޡ���w�#���|�r��u���E�ś>�a���w���SN���9����w��Eߏ������7ID��}�G�Z\3�,��֍g�P�<k�%�a��w tӏq-gٟ;{���t'|Е���$�=���<�I��j��I�H=�L%���kRp�mt7u�z��'�v�*��ή
�}ɉS�~����.�s�ɗ�r3���!ڲ߽c��/�/�˨@�δ�S��^W�9����;�r�c��O{��{�^	1�p�7z����U����3�Eѽ���O�q���=�y��@E���wj��Cnj`�(����ꢫ�Hb"���<ǲ�75q�r�
���g��>��V����܎����H�/�ciC��u���\[]�c��m���ɡ���<Z�5^4�7��$��1�[��w����#��E��o�-�K��K����r.
<�Mm�ܛ��._�(��;�FAqnj�eL����cR���o�D�l����jc,Qo�G'��^���K#f�'��8���+�"\�㑸b����'IӘ� �C�M@d��G5IW��[դIJ���eG,����c�IS���-�a��0뇔r�/�#\>4�G���ZƲ���DX�����U�ҰGI����9Vv��tk�sլ&��F��6����,}�Ԥ�v���3�P�>��KM� �������7����b�����υ��D�|p�~���w�������n���mH����
ՁS3D摦��Ű�`}[�����gD�~���8� �*�Dm��@���Qb|F��i���Nh��눵s�Eă�a�d'���%��Ko�u��\�V�:}yY��\`�LQ����-8a�e�a7
MĻb6�J��
b�b�����	R�AƁ���ɪ�P�xt4�A��!�n��Mb��(�Uv�T��%�[�	g�7W���چ�ꜛZXL.>x�߱}�yŕ��Fw����v��[ov���ٻ�-A,񴅭O�*7� ~�অc)�ul'}G�,�3ȃ�i������u�A8%�6,�&�I�Q7���J��9���2+��/Nκ��I���֯&��?p�RB>�{��W��k�K��MN��;o���w�[�YM&Μ�(�w�C���d|���������'?5ٽs��ӟ��^v7������Ç�d�,�SG������466��o���<�9�XP���1�<���;q�GU� 2N�_��7���w&Ǿ���/x!kC��?>�|��_2���j�|t%�\?��
(�YZi���&/�D��W!���H~��:D`í�����N�8r�+�/������������*�{��K������=��7���q��>9v옽��ˆ��F�	K��֚p�����woǟ�����M?��ɛ�{R������s��z���������=|����"���h������}G=Cds�PD�A/�ފ�*��"Q��
rF3I��	7{{����q'(ԍ���,�/C��{*I�R�u�7ip�D�8�Q{n��������v%Y��AF�0Ǽ_��H^�s����Drn��>�Q׏>���r{��}��1��z�u�/�����n��T���:f��İ���4BN��:�y�̢��Ib�������Z�V?'��B)u� �݂�=��ь��-3�q�;#���ì�
���2
�f9�&;�a��pDbnK-�v5<i"H�@h̭ZUJ�^>�(L&��~�33�V<l�lqI�>�enM�v�1���Iߪe ��^���s�U��zْ��� ��dHR� ���g�����s������2B����Ctky���04꯲��e�LR�0� w�B��/�� ����(a�Z�Y�̒��{O��Z��d	�k�=>���b�P��_�.F������C-0�y�o�����%+N(g������E�E����JNeR�i��Q���B>[?��4]���P���3�$3��>��2*(�+m�����e�d\# ���}e1�F�!/U0�k�2�{��}���R��ὨΨ8<V� ��=�����3��)	/h��Za�FI�V2Bz�S��	:f�.Uk�҂�?��� �70}�Gz"H��Ym��n C��:Y�J���g�����$�3��^�Fj3����78^�'}�@�:~���\c��h��R�5��W]9thr��k�ܮZ�H��fD)���.�eG7�_ZXt}=et���G�skp����hh��7���x���'��3\��JQ��`�߽�m�Tnj��r���XH3����ї�N�Aۥ��gxF�n��Ԕ{ӛ����O��7�QЈ������k	G3�_�\r����}����d�Q��A}���LX.�2^������9VC�v�������^��g�#�42<�v���?�WoG-�oR���_x��ϋSԑ���J���B\�}����54��B�C�t�� ����`�%Ά���p��E_� Ӭ�>�B���0�E�k�!�=��v���C��Q�&��n���ғ��Fz/OG�:��)��"��u���s�����}��n.��f#c;�$�JՁ���q�]=���F�/������F��x��;!P�ܾѽ^��aA�qhO���{����[_\r'�?|͵�����/,!Ԏ|/�
1�v~�m.�����7k<<<��uu`�֫p��n��p� ��K}N��r_�ua�!w�'y���8>N�$��ii�2��pƿ�g~��7:ݞ#OH.����~�-ɯ���
E�u���TK"��I��n��-�Y��u�ω&��Vk�0Τ���25�-+qJjwG�t�1�<��#L�y��|��]����5}�}�F@j�tg��Vd�����L�j�e#��hL�2aКƩ8~��w���hʙ�k%�⑇̥�X���1^4/&\y�g��JӞ�j�_����F�Ra�'��y����c��<Z,�s��F�aj��~ޞ�ؒ~Ĭ.,;�?5Cʶ(�9UXJ"�t�����t��y���S��V��c�ѼT������q�ԝ��A��� ������c"E醶�D4^i^ ����
��F���P���N1P`��TDi�J�o���M�ET��#�ƛ���+|�� �Y�-R<�`�,鳓\#f�޹c����9n�4yu�G"9�qkIG<���x����1�ՠ"��t�F;R���y�P�h|P��\+�;Ú0�uaU5aS��eg�T2�r6t�P�r�9(h0�k���i��9�1��5w���I�G]�u=�8�'�<���������̸�TFe��O���z�K���m^+�=>��-KWu.��R��� R���=��Pƻ��y2n���� �x�D�!��C,�\��_e8$C�Us}����uW5�?Q���э6솻p�2۽���#�p��۝=q>ٶ�ɓ��Z�e�F��O}�3��O=��񘗆l��r̔�<}�,�:�+���h��:t�	צ011�8�\���t,n��z�W������9����g���]��/~:y�s����>�����%�:qa�q���|er�=oA�%A{��_�h�M*q�D,B��/
������i�I����y��N2���~�i|�����n�F�>����~�2���U�dzz��v�m�j������FǈG&W%S���cB^��)��U��Y۬����Jn��>��~�rn�Q���n|��A�&:�������G�^MF�������af��?�Ӝ��7�~�7�&����مY�9ʆ�م����,��
;ys������N�2��y�un�1w�]��1:WFf�z�7��ߒ"O_C���+u4���2ʼ��g>�)�t�A��C��N;�,��M�~���S����{T87�x/oB�S�!z_d/Eo�B�N�4&�Ub�!�l��:6A�68�;�ˏ�-���2�E3�]ʌ��L�����iw�O_�+��`��H$A Y��T4��3\D�$�������F�)�jS�M�[��Z*'�+���i�P��x�L���w�>�=�'Ƌf�f�ҌK�=2�l�3��D{O�f�jU��Ű薹5}[�Ա��m���?����1�1�h�0kԬIcz[�7�P��-��O�o�Ȋ���vU-�01�2)BF3���P.�ǂf��2��R��i��k
��<�-��V��S�VX��+Y���=����4R�F�?�+1�j��=���ZuJ�"����0i0q\���Pa$BC��<�B�W��C�oڊ��U�7�gVW�:/��w `7����&�4@)A�� ��+��tyq>��8i	���={�&̰�8t�I���=��T:��^7aj�z�2u�\��هv�F����Z=<��8/�`��5�"V.�6qd��S���x��������{��u�w��L�}F3�ьF]r\��cx!	)�����	�)�CX`�7/�@H�H$`.�lc�ƶd˒�5#M���L�����=�\=��n�y�4Ϲ��~��_�2�R��|N�� ���P�]�Q#��j�$. ���l�y�۰q�{�ч����1������9|���Zf�H��0�FH�4�?�1A&�v?�c�˰����Ht"�L�B3L��$5d���0l�x05�Xp��H����c���~�����ɓ'����q��؏!�.��%W\�΀}�UzłU04c���o�K�w�����	��dY�d�P�󨭫p����0X�i�+�l���	m֓E�'  f}�Vt��0�*-��@�S����Zﯻ�j�M~�g_��r���g���v_�����~�͌q.Y���>YI���B)dy}��p�W�䨆wk]GՈ�/�Mc9�lM`{����a�ς�i��x�m?����V���R?p��=�w�S�������ݮ���O�պ�������&��$Q,)�<aȄAc���;M4�jr�hu�K�����w�f ��������߽߷�/wӈ˓���nt[wl��߹�bj���jC�ʤ��bP �I�u��z雚�qgN�L[ �DY�s.71\$ޭ��t|?<c�7�ݷ���r����u�l�>�|L�]K}���֗��ҏ;(`^:p��~`��}��{���F߹aS2r���h �	�fq���}�NА��Ѐr���"ȸI���W�1�R&�4���i�������@T,�R�L����=������DW�zb��~�7ō��C̵ߘO6m�/��nL��o��<b����mxPA*I|�*F������%шՒ�3��Kf,����lܡ_�����/����}/Ld�Z���_��ҾP^uTa�J��Ʊ�+̎�z���=i~7ػ�+_����e�~�1K3��>�|���K1��n��-�� �ރ�����Isջ�艮޳��}�'/��]K���ѻ�]�e���yO���͂��e��<�1��%xRjv��(~t5���yAmҪ�a�7~RW!!1^��w���e,0����4����@��_�d	$# *lmo(�c��s3�YL»=>νs~#�KvX��Dҭ�bs�c�il�40��`+���YLO1�!K�3��Z^�
�gvVa- �����@�AU�5P=�%�F1tб�������b�6�}�&�, ����.��!��7S	�N��o�D* .A��q[���g��f�\C��U0��w�Ԁ۸�-�9�˜r7�x%�CO�������:�Y�bOK"�� pOem[@�kN=XQe�]'X�$Vc�댯oXGVea�7��z��~�-�P��{r�^���%�0��<�ԽE����u^��K7l�w	�A�M���GE-��
$�Y��S9W�D���,�]F��m����Gl�2�;�x }E��rW^y�;|��)�ܴi�$��y��;]�m�K9�5��������K^������r��뮻�w���^��[�-�:QD�rTNc���?��$�L&Y �`��r����Z���w��n���օb	R�h�A}
@���ʿ�O~�R9w��!w��#�7�������`�fO'�����w��sWR_�L����T?X�wj�4��U~۶m�B���������?�=�� ��_����n��B��=��w����������ۋ.ަ�D��DU�aJGЭ�\
	��=Ws��>���2�9�"љ��Мk�)s� ����.���vnB�`驅�䲋6���*�б��j_	/��+.r>��$\3�xo���VuS@�GA��h�I*.ru̳ѡA70<�k�7K� �"H�C~ۆ ���Ձ��a`xŘg��,����W�atk�˪X�m@}vٲc�f]D�ȗ�h{[|����&W�z���'�F���b1^�w6^|�n�ݘG,'~G7�+~6!��3� !�4��! I��U.�E�p�]T�׹p�Bo!�I��l�HQz@�ӡVX���f�Y߅n>r��|qb~1<&)���1���p�9�#� ;�b����RW3G������C.	�(��A+?SHL��X�:��:1nX}ԍЇW`C7AD$Dv�M8j��.)�w̋XV�}+O������a"�dߍ&�"�B�w�����*�Tiz.>��RGn.�X ���gnmY+�*b�k~!����Y��U�qhc�uUq�������b��sۑ�b���[������OK!�rP�0�.L�jO9"I��FF��b����[iZy06i�����h` ��k})�n�ʎ$�L�W\�#��÷Z��W�UK.����Y���G��/`�8�����tZ��!$y������dtd��4���@ʝ��%�p��eǋ�@�`��g󗩉J��Ul}	� Qo��ⷐ&$��ص3�GK5;Mf%j��|CmB1�X�q$�'&�I�"�l�":��8��1��
���d7`x�º���}�S���O:�e|V[Y9|AK�V�ɡ-��ʕW��	n��I��hUw���\��I��
�� ��|�}Ly֢NB��f�Mt\Xv�"��� Ƃ�
;���az�x��@�,'hE@V���½��G����o&��/��\r�ͯ����d�ŗ�����Щ���g��#�ƫ�$���/��}�����aY��H��_iM���?68��<�WV�y�0�"X~&0W��	ltRG�i�V21:��T?H�M*�>3�b����&����߻w����b����o��U	�	_�d.ٺ�> �J����B��&!����B����vy� ���K�A�S#�t��`�*���a�׊�f��A��θ�[[�-=�Gڛ�{���+^�j��Oݶ����,l���?	�����}ዟKzPy��w��L���k_���������W]���!������oGc�����6�d����S�^��W�9iM���nw����䟿~����j�}p|vŵ��g�H"n�����Ș?q	6��r�O&0_W	��|�ddl#��O���|I򮷽�w��L��G��'����8� ��I��v�O��3��*�6�p��Ʌ^��Ws�;源@l ��ͭɖ�=���[��M=���2�@Ŀ�5� Ka4��E�5��`|�ɑ�c����d���2ϊb��7��2f.S\���u/�%Syf��[�"�]k��/�Y�s��4�Jw��//���q���nL��S�n�6m�$��l~ۋ�%��M��l=��S�2�x&��`�J(��'_F�U~&ѹ�c�L���g<�x1ι�QV��i2E�_*��e4젴cZ�`̏�4o�|�2�:����~�/OD?XP �C�xm0x�	>�h�p����R����\��e�V~�Ng��VGյ0L��!OjKnΰ:�hrδi��S/���Ԋ���e��1����'E�?c�g���W}�\��g��')�c�O+ʑ蟐w
��8ھ�6\B �,[ kR�N�%�Pj��b(E=
gA�K,�	�幙	���>�
�e�Z� Aku��!!!��"�a-{h������(6�:�00��X˸HC7�k`A7٪j�\Bàp�@TK�$Ls �([� L�*���ժ���A`�d3��:)�/��zA&􀤃T_2��{�ZZ��P�C�_LmE���+mRSW뇤2J�)�
<D��6�Ҍ]�K#�_�1m��D�S���i�{��%>-��:3��p�z���Y�$\����o'7�����u=�/��M�CG������F0_K������hF'�� ��X;11(
%�d="㌭X�!��8�i@�:  @ IDAT`�ϳnso{r��~x�)��Q���¤ @�����=IF�C��S+���� @�&���5 ���o�������Q�w�����xY�	�;x���YU�����;�Zi���"ͩ��j��?�wAZ���>�$�Ӄ���b��$�y���w��M�X��x�vd�c�Ӂ�'��$����fEkk+Fn�b���ر#��{�v�����9u��/�~�����dN�$�h�H��e�5�� xQ�	 ?39�kQ�8�v����e��P@
�	VR�0r' ������Y^p�[���<�k��e�y�KX%�"�j��q4k'��|���p�(��'`�t�����lnpM�����o�df�m�hB��i�2=��{�I����6]�hO��g��E{��7���v]�7m���iǕ/{�k"?)�ݾ��� �rho�������V_T��ɻo�s�x`c�Rȡ��7���	�a�.7;[cZ�,^��ɾk����{����D�sō~r/���1m��w6,��F7��0]��VB�������j����+�ZZ�����֞ŭX79- �a��.a���r�f�b�f���
��r��ʫ��q����q7���8d��[-קθ�d��č�!��(}�{}|�Ω�o�L�w*��*� �O�8��O�U�����ӌ�?�E{B��NyrLa�4�v�Pmt$�����1�|ޚt�9w���t�~��AP�k��Z����pf.;O>-5iS�"cB��8z�.FA�Cy[}� 'b�!P�H�ںº<���#�c��3���0�m��P����!�@�7�D����Ĉ�Zk��3�I�����aNf�)9p�op`�.� }������〧��P� 	3`m�Ԇv
@�d$�5pP,\�r�p�d���*�$�&Fa�P?��z���F,&/Ġ�!�	?&C�0�.IzIID�m�K+�i�&/����:Z�k��C7r���Tp�v���4��C�z�* ���w�0n:�c��r��<wп��/3"i=0�:8Ef���"���_t���TFl���8��I��L��� F,d�]t���Ɲݹ���܎]�������7��޳��ˮ���~ֵb|�����s�����=�U7��>���]�)�\�:��U5�Dc4�j0t� 3zù����r*�S��������qV�^����_N;W�@-���>��Ot�"�6�,.��׽��m��Ss����;�.�����n{�&d�:��*e��؀��0 j|��Z|-���!rߙ4�6�g�~��wop�]tsp�Ϣtq{MeM26f���:��|���A��3N��o�q76�6�͛73_*������]����T�n���/���������o��۫n}����ˏ�&����,P�J�{�C�+����� ŉo��1�R�0=��0 o�0������Z�?7���	����������|e34Fz�$W#�X�V$�а����!^��������M�\wǆdr|��\B�j?<p2:���	w�Ghj�4W�oσ�����O���#詪�6�f�ɻ�$�-k�3O>�>H?�o��]w�I=&IsؓC�BݺFׄ�����Tq����>�JQF�e�=����'�0�BU����v��.7���'�죴1,�~+��bx6}�?W�&W�t�=�g|�q��ha�?&����w���D���`�M�6=�%&���A�f��@��Gr}���?V��ߒ�'�_������*]6m������o��Q����zZ�tsM�*|3��gyM��G���"ML6��b�c���i�� 9�r��JRdg�����P
�\ic��m�+�Uh p��\ ���(?�V�&�~V����*��}��E�=�i��[��J?,�0�c\�ʦ�=�E�P�4�&n�~EYS��u��4N��*�v���/��C���Y����L ]���fʲJ�2b��d���.�v��	br����vf�+�> �ڎQL'���X���Ш@$� ?��~����+����+�H��@`�1yJԔ%w�,��"�ʃ���`V.��X��@h��S0���
�>23�<A��N�&�akț�W� ��*�$ǖW���"ю�`|05�5��RGt�7ɍ7�����[7'�[����մ���:~	Fߖ��8�j�� hBJ�� O�!Ѕ��xĊ��-�pn��U��ר��Z��V��N/BB�L<���GK���IwՋ�&���/����7�=���6m��j�������O|�]��1+b0w�#�]9��9L�T�djb
�P%��T��ȡ�q�Q�p��%M�ҪitM@j+�����A�7d�_@z���&'қ��5y���E]$i8���'K���l���ܡY �^�03��$��۷�HN�.�����)�/���j�4�Q5�ºnuoX��N�΀�n����4a_{ݍ����vw�y�k|�(ـk ��/��׹щ9�<�/���>�!���{����7��Ͱ��%��������;i�f^	)��|��!�5 ɷ���l����9wr��wu�b�l�{r�1��/|��?| ����	L����IK�ySw�$
>Ň�Ocsv�&a���u�l�/$���)��2-3��z��55���O�����\����O�S��˯t7\w�;|䀟���-���t�?��Y���e7$O=�C�e�&WQ]��>�7��W�r++nC��Io�]Œ�}���g�J��� �V�_��7%�HY2}�P�	�/�>W0A1�ɵ��L��y͢s�S,���m=h_�_�H���w�=��=�S�6��n�W�J�)<���=ד͋݊n0�Zh��B�˴�usԣN�MlC(Ïf��L�ӟ���Gt��������������}��_t��̷}r��2���l9x3��/_W������0=VN��Il���W�!��}�v&Eq�q����z�ޠ|d��q2yy���F�Jc��!��	\"�����n|rE,�ʄ��U0̢\1Ze�>�����,L�O��d�_��i�♟p����:p����q׀	���[ �3~1�bi+%k���Z ��Ny�vX�iޡ=��v���Z,a���[Vt(?�wj�Cݶ�M<d'�K�O�ְ5Yi�XXfV��]�@�@��"E��6v����N����k�!���;Q��Bs]�ۺ�׵c������7��p��)������������
�s�KP��`�M\�x6[����0 KH���*_Y��NY�W�Ѻ
��J��V�[[� )���&
�BH�0��T扸0�
��K�7`��8�L��"@L�Q���2M���>�'1�z�ˮsT�i(�L�5- ��_�˱��:��P��W���1X�w	�ԣ�%�$lz��8��x��iJ5�Ԣ�`�������}��?y�!�]�:�?}��\m�r2z�9��7��|g�z񅹶�.�Z	���1��z"��mך`�kQDIt0U�$��¤�$��C
v(�* �tvuA��L�1g��T�_�b488�dX3�;����C��Nu�|*q\��I����B�i�B����<MU n�Oa����P}Z�6n�(�|�t*"*��̀=�J*�r�#�6>1�4��̠��y�w�u,W׵��<�l�~��羇ܡ�}�I�R][��_v��_}���oq�<{ rv�``��w�v� <Ã��y�Y�L:����H�-��.���5��]�\�ͻ��Ӈ��H?�"�����a��ާݳ�@�~h>;�w`�ȁ}��t��KDc�0X�F׼U��b�c�M��A���|3@�vw�K��������^y�������?$��A0C��%]{õ�@hw�39�L^z��n�o&��+^宿���L#�Y�{7����=w����f�/a���v����w�_
�����o��{NL�H��!��J�SQB#����܀H�@]��1gv�m[�����v��_�.�w>/1޿�/�),C�1�°K�%�T�3i�C��G~�.Wk��ȉGD�����2G������/��ξ�W������G��Y�lX��\e����j�6P�}g}��푟����a�jd��v�3i3�˶�&E� �'�b�������Ɏ��RQ�W�˪��Bb�� ���BB��sY�2̖�I�/+�E�kee�f߳�c:�#m��.���DjQ��Rr6�~g�,��9;���e�7+8�VX��UW�*,O^�8���q��-{eg����h�ų��6��P������7�Â�I��+�4Q}`6f��R�|�Wـ�Ϻ�$7��g�b(j�_��`����3y�\�a *U^6���V�ט4� �0M�a����x�,�AH]��l1��|�6%7L�'�5���\�Q���p��Z>¾�%-�I�A�[�a� `�""�op�G��e��/���z�#�!�.�:���Ϝ:m��(�pX,LT�zm��4-����#�^���bcBy�4�/����G�4i�� z�x%D��`�S���ӟ��������[n���ɏ|���[��{�R5@�.HR9��іiPC� N�1���@��S�H-U�%hkā)�6�0�1��6cr����S��Vi�Ȟ��&`UR�f�!���ܶ-��ѣGm<&�	����cǎ9��?x�یgk��?��7`u��������X��VL��fI@�
@��� խtS̩������l~^���vS�Q��r��G�b�ab.��
lM��Z������?LN���oy�o�i�*��dh��/G���M��I��94��˿�k���K �"��Ow��~���)��M�v�G�!O�o������ϻ��i�]��[:ݑ�Km�_߲͵�pI`d몘�#���O@��v����Z�Q�9*��5w��Qx���Q*.�Ln{�k����g0:�̖߃�ȵ4���^�j�����!̄,�����_�s�w���w�y�H�~F��rHc���#�N�Ɔf̡Ժ�~��$���y�׹���[�FuϞǒu����|�K��ٜ@f�:����-���9,�,��1��&(���d,+˥��ɴ><Z�<��>gO���0�~���nL���}�~g�,��S�����U�Hn�����"�u��%R��4x��$q���Dd1�U6,����^�K�䡰�'��k��գٰ�_6,��8�)L+��ݬ���_�Z�V�l��wŉO��:�f�@��V'�8g���%�-���Å�|�lwT+��D-y���m�{�3�M4�`E���ߪ�J���3�E������'�Q�6�eܱ�	L1��`y���ˆe��n��xY��-me�t��xԵ����y�F���3�Ud�\h�Ԩ£C���`��>%���_YU'�|��V>�ȸ��>�rA�9,���b���d�D3����B��K�
d}� ���C���m�����F��`�6�UDߙj� ������m�C�j�a�#_�RN-���h��K���UW,H�"�D�@?,�"F�$6pA�����B�<S�5%�HN>��"x�CX��ٰ��T]2T�'}K"��Fu��G�������CNͭ[���!�E�ʪ+V�0��?=g��qB��MQ�ʲx�VQH�JtIuAIqER�"�Ð	`�+�H�ꓰ�i��W��T�vi]x �"�AqSs�u�Ec��?���3�����Ƌݗ?�)��/}�] �M�^�1��`+�⮪�>�r��;4X8 �1��ѭ3x�m�!�b�V�����T�c�=]X�jj���A�ZE��Ha�_~sr��o~�b����7�6��&�����v�P�{���毿�j{�6$�RI`q�<����(�YN���΂��j|K�i�5ԯ"<P��i�Z�aڡ�8����a����%��3I'�2����=O��'�>�d_�@�6L�`����;����_~ӝ<~̀d������_u�50`��x�{������7�=��}�u�s�͸�f6�*�Ѫ�Ɂ�d�Ȑ_��jw�/XA�5� �D��F�&N�s�6� p���8�bh�7�3
a	��~/b��+`
���Z���gd���t����������/���cM�O�q�?�<�o�ookC�A���{�q���B�I����`ۉ�@=�w�k������S���Ν�����-��OaN���ւ?�tdt�m^��US\TUY�fKʓ�b̩ 
�fAz�t�!@�,N���no	�6E��q��V��G~�Ed�
����{�+���+�s�����>�Ʋ��&	.[ڰ������P*CR%|+
���ҍ̼����w%��(��Î��s?��'�����E�1?��-�A�cU�������NW���ؘ��E<K�I������_��,��|���a�SaV>���.��cǼ�p
f�ƭ�a$4�'���r�
���|E�>lp��I��R��K��*`R������~� d��u�X�,�dˊ��=g��\��d�5����i�X?e�d��;_\�"��ajd�3a7��QdF\>z�S}��;&dHVE��s%� F�����~P�@  ��3l��Q�
�	b��H�V�!d�� 
^m��(�f�D&��6^��e�0A4� ��T��Bl�tj4�X�"����.Q��7BӴ��Xin,IK4��[�"7�a�CRW���:����H6m��f�l�����Fl����'?�Ќ��f��`8��0�4s+��A^ 䨲q��6_m.�e�
ռ�����?�p�i(x��ɪ*�ڀW��3�{p��Ϲ�~�o�5Wos/������\w����w�����7��'5t�����k��g�}��{�Ǝ���� _�,���5W���6w׷�����nM����� �V_�Z ��0w��(��R_{�J �&l���������7����6=O��s��䒋`�YF����	�:3��yt��J �R�YR���mrÓ3����]3��|�C:F��W0jW��6��L�0J���(t)$�:@}F�/��W�5�+�|��CZMؾ��qH����?���o�#����
4�� J;/��R��o|˽�5�O���g�%������[�k�f!?V�e{
,�x���\���$ݱ����-�y�.)�i� ���Q �rHv¤��FW׶�u�G��7>�V0:��ZBj������بm]���..��Ԫ(��O|��1��57\/��9t���r��NXоg�q����1ӌ�s�N������a�f�˶⁧��y�}
 	,����;!�v�/�&�o&�={���ys�c�V��g��Kw�� ��P;�i�R0S���F`0�Ά��at%��Mr�D-�0���c���p�ˍaz/|b���c�l~1N֍��_�W6]|מ��;�.�qe�a�H��l��͔�Ԗ�vt�������������\6d�z�P�^�K%��)cΏ��.x��&a�7wK�7�9+.�o��Q~�𘿹
(xbxH7��S�S���u
��rh��6A������8~�SZU�cӉB9.��ŐY�$'�=�.{0B�r�Y4P���F�:VE������-��USd}S1}��P?��Ҥ��G_�����U�5�_��P� c� W�y��`|�с�Վ�h9�|��z�5�r���kȝд��U��o�./X��VMVj�Sb"��hx�q���P���eVV;;���o1�	�e�6+�)��)�v~ɘj��B�UJ��e2�f��|8^����ыS��h�j�� #qp����Y�f�hQiy�2����q<��X�˵ޤ�:��9�whT1|k=�����X�3mR�0�2��e�'�P ?�c��N���?���X���2t���X��ol�����:3ZJ��z��f��"ѐ����ڨ�3���D��t�d�`F�@;#C��(i(��l "������PS� ����#Zm���1hv^Ԝg��2`��z��K4�@�BGy��@��5��ŽޕC�X��c���g��!���C>����^",���f�H<U`����pHL��Q|�_����Q���=`ĸ-�
a�+Fc8g�l0](��Z���-|(!a��[��c�*���B)_��ܽϸ]�����+�{�{��+���Ns���&�yן�ђ��F �r��?}������.w#ë�}M/M���'m��-�����w�~@J������Ϣ�|CqUr���oN����
��蔌Q��}�I*Y�O?�Ϸ6��W�����><�.S���5+�M��Y���K]}�E���)�G��6�'،V�+�'�Jz��1�{��\I6Bn:��q4�ϛ�T	J��Ix��I��P�9C��v�h��Z��|��u/����ML�bSx@��:��jmu]�QL�p��N�&$�fF� N'7^}��1�U��I��N߅u��rhHگ�o�ns�M���ze��_0-���L!%�͟s�=�����k�h�jr�̤?6�qު��6�! ��2��+e\�U6gc?:��ߊX�Ip�'�����*4�����.7��T�)�2��7�����k�u���QS���)$
���0�S�*����'�U5~lXj*W����FGؚ���h�	��ڲXX�͵�$���3�uy�O?�����^3�����r3�%�[Q����_V#;��V��1�k�_a�?u��hy��
>� ��z�պ�Q�l��wtC������̆E���K�b~�?��ͧ0�0,�#�V��>��5����B�$��6/ޥC-�DaXQM��>�_�\kX�@�;�G7Fa�?/͹�b��f�9߻�ưB7�s�����GW�a}�)CaV�9�~|�tz
\Y�0h"S��tƨ =�.�ϯح�ܔ� "��r��zb=b��۪�C�i  $1��rC+�_��s�_eQ��U�5�C�VP�1�_��'WU�~�K�<�|����+�*1݊W��i����)���'@�p2���@C�*�
�:���:�y}b�VO�{x�s�8VƁ\�(��<�q� $���$�&X��#���ɻ/Č��+^ �_�[@��|eaI#�k��[x#�&%�K�Kh|�򃞫Z��W�t�;3h��#	��~	�n�$�,Z��2Þ@�r�V����
�Ecv���<�o���@ g��2�Gl��rNb"iN�Ա�!Д�����Am����
��t��[��������`����{ �e��K��,�,�EZ^�Ys��sɋ/�ؘ���wu�X�G:��F�(�2��{K�hy��q|�s2"�n�q�͐šjZ��_|rE"&��C�m�0D�
V�`(v���?��Wq�7v%#X���Y���&��t���~_ �� @����q���!yS,5`�$��e�V�o����{����`��G��'�tw�u��^������֝�����z�\�u`6o�q۷l����*$�D.Sz$��d�����=q��s��o�pãhh�)�è='3 Ma:sA�tn;z�ȷa���Q��:L���Y�1U���$�S=�8�����:7:=�5��Y�)�L�{
�ni������1���t� [5����|�?��î��WX/�ַ�Չ�$@�]�z�������!s�I"��c���"$�'��ۀw�y����[S�I����w��~�7~W-��uo�_��c?�0A��9װ��@!cY`F��੥-��Ј�m=J6l��f��F��5�Z�t�?��Û��^���W�"u�rY��q�U���T&P�v �p_��	���M%���%�)��4��j�i�
�R��@��k�[���4�w�v�����.nݘ�q��Y����iqᣭIӞa�˨rg�X����ģ����]O�wܯ�_R�_�Ÿ�=_�Ǽ��*��qye�Ÿ���w�uHEAaSC�B�u0�XnLՆ�c�YT_S
|��@ �"b�a��_馿�IO�&���up��%W�o��H�*N6���i~�wL�V>[�er��ˏ�ou�P�$����F��"�>ƌ����Ky��t��I'El�}g�QK��O��Ʊ�,Tg"qtDcYE�U��m}Yr)�j$]��j�lA�ǎ2Wa�D��}g�Q��,���I�R�Q1�A.Z��&DG��U�ű�I$��%*_���V����=�,_P�MhZA��iBĐ ��H595�jf�j�q���	4L�d�bÜ��e���N�B����l���F6��ZGaJ�BUQ���*l}E��"����@��Zn?!��VH@X+��yHW^ra����x,�%H	�S�V�~C��(Ҟ@�I��@�	P�zt��x ��)��l���j>�4ګ�T���5�(G�Xk�v��v��?<:C�f�U�K܁k
�?����O�-� ��q
[E��Cf�H��b��iD���d�Cp�9;�-E!��p����ǎ���C��(Bd\��A��m��(H��jz�� ��z��V����
�U3��"��������/���Q_�|���'��%,"�����!{54�%�≢���P��\�����G�k_u=H�Ugjks{�=O��Uo�����:xS��y�����FΌ%s��8z���[ts��Z��y-F���zuzv�������-�/���x_j|�;����lg� ��ˡ�2s�RRX�����6?L�����a�'�H�75��eL� p�Ο�]���Ĝ����\�?5\�cG�&����H&�q���핗��aBF����=�{��|�����d�ƍh�_4��3	����$M?�u�]�h3�c�����Б�hʞr?�`�����,���կ��݇����'�K.�����{z�~����x�Ĕ��Ź�1�73Wโ�,gdf��ü6��SVW�xbƌO{��0H�xuΎh5a����?$r�䈯`�~HJkC�P�z���� �����a���l��6n6�a} ��}����n���.z�İ%<�:4�f�nV��v�I���Լ�Gۙ�]�պ�-Y�1޹ܘFaٸ1��&�J�Ҹ��hǂ�Ӗ� �u�����*���(0=��$]�W��>1��s��0�ٸ@*��w��\a���d�<�_�~�q�*�b9(�=����Y��]'����V>;��ӄ�����Q�h�9]�.�(^d�����b�Wg�W�e$�(,���N�|Ni\݃1RY$�����9}5��n���c`� �_=�ZU,�����*�bX+�M�e���L�T]�Zֵ�7���n	Z{MW�<�9<�M?�N�,kk藈��p֥�!���"K |��C�	$k�f��L�"�%B͛��HK��9���H#�MaV��:��o����&���y�/F��h
�W)@�<D*�퍑f�����o���~b����}ɣY��3�L�2��i��C�?K��E�A��g���C$�D��~`Z�c#�3���	�|i6]�[Q��m`@@���W|-܄�N|����{�$�k���OZ��_� �Ŵo�V==�hxuu�c����E���*$���С#Ƈ��٥���2�
��U�u��-�%��Bd6tK�fPHiI�k�Zg����QT��W�p8rJ��(yȶ�k*в��MÐ\
OJ�L�9���⊢U4g7����pɏ�g$��)�W�ܔ,�#Ώ�b=X�o�4����sF���-%��k����.�i�&'R��HW�D��G��YEGP5X�u@���9���� %.c+������K�ތaT�08r&�oﱳ2c0�J3+��Z�t�n��B�p6��2�Z���Ḱ��ں�/�7 @-�|�M=�`�9ȿ� �Q� >����A�K��%�R�,
sh���� Q4��@ ����=u��W��\9�p5�̐e�xv&�«E�m# �4��w�.܆^�7�w�}�k_s?��6�A�e�T!����F�K[�mu� �
Y��'c}H���d}�F/~��-�h�.Qm���7�,n,���~�޶Ο��3���眑���M_�ր\Èi��񽽽��_n�)��)���A_�O,�US�)}X r���0�ĥ�񸶰��"���z�l��"��ҡ5�Z�&�v�7,�P���U0���6������f���G��]�+L���S�/� P�*��:�`��C���^CS!�5�w�gmݪ����aTiW-�1�k�p�8�[��y��w,�?�|�kuvmlC���ӯ�-�s^tԣ|�X�0��K������Jf<K��xY��d
9�����iv[P�p��eErb�� �@u�$@󠁥�|,R���S�>B=�d�u"���x����OOk��Q2s�y��]M��!h�؋Z�y7�x�6�Q啖k�����-*�s�OT�ꑺ�Yâ'��l�a)"CAZ���������]������8��]�����#E����� /��h�c�&�:~j:�Vi%�j�,|�6lk�K�I�Vzb;B��	�ުe����{Y�C#� V⛫�Y�A��k~n�[~�I?R�Q������Օ�$b�0ߦ:)#ޔ;C��G%�ʫ���NH��2�MI���Z���/�<�e0a"r8�����(Ռ�"'<"�Qg�dHZ)V�CҨ�t�$e��A���%k|u�?~��1��@_XBELR$I*xR�Wt�U���7���)�!�`G��B0�P�����1��]fl-2ڌmF�*��X�h#IhH��IMy�j	����Q�<����$d��#0��ψ{ף/in�;�cRR��6n�dڝ%���	�����ػ����?�zꩤ��۝(h_����L�$Y#;e6cBu��X��bNk�#���YT����j��;����`̮t�c9� �3U���lΈ+U2�e��	Vi3*�`�_b�q��&�O���)-B7ubh����wv`�?�C ��d`��k��d�k!^��nt?���*cT>ї��]׆�L�%cvf�Iݗ ��?~��M�x����<7?�J�v/}���_��uw��[�F]�~�~��t�U [��U�͜r������:��}��
�D� d\B��R�Y�}G�|I�BU����9�\,-a�1o$(u��1җ����˂���	���_�O�^R{"��$�H�"ﵴ4�r)�t
�9(�D�U�� ��am0...�Z$!��"�/0�%Uj�D֔Xt�3�����rp"M�6i_�{|�N�E�w�/�Dyd��2�
�,#��+}���i�Ș���\����?Z(��ne�t�­P<ą�\��)"O�(5*��0k�^���c���{���?�|�_�EG�v���7�z����L��30e�P��;��S��Va�P�p��'dĕ�Y�[t~2O&\㟝�Fa^ʁ-fD�p�A��`"ٳ�C~��2_>y��u�/T�L�!nZW��x�%��,]SV(��ؑZa#Bi!�L��p��kRQ^�ͥ������ٸ�-�����Q���P^����d�P-�nU�V�4�X}⵭�`[c^qc��jIAh#!uP�功��O��*ƒ���[�W�/R*(|*��Q�$|�F�!J
�"I��|'��u-~��s�(p�>؎J$�^ ��e�� �X�D�`�0W9��vp��_`.��|/N�(J�p��=.�j{�"jc�����#:�d��G��H �OU6,���E�D'�R�� ,�u!��8�X����mo��v�)!i������?��8 �M�ԋ���%}9�dR�Z9���L��qY�����OL�"Y�?�	&��i�S��oƿ�id}f`7C�O�S�&3�M���2������샭��a>�r�Qҭ�D]��&�	�4��8�� 仫7�aJ��_�_�4�4n��>��<���ˏ��o�h��h�{R�3�<�r�N'x��w��Z9�u�#��[��@� E���̜��iT����X����$`��׈�Cr�E,J
?K!�/�t̢� �/��������n���F�Zxa�@�P���И�VI��C��z��}`���z��M����vH}u��V�u7�b����	�uw�}]<OuLP"�)`�������KK~^�=�zzz�#�A�})@���C����B�N.��w��A�ۻ�_��������#?r�ݲ��zX�MP��6�8�j[Zů�L"�WV�� ��xY0&���i�0�-�HP2���W�6$ޤ�J�0���u7�%3�ib =dBa�4���^c��Z�\Լ���όyM�.�;���4�3/r�_./�1,R�n��Ӛ�=`��"�T��CH���Z䟔�jl��E�v�~ *e�)/�������JЏb������{�_�����_(n�q���O�Y}�'�׷�QEQ��yPq9u<�XI�I�0����S/�hz�<yc��{��4��+���I�q�zb<yڦ��f���(��xэa���zf�/���lxL�e�ԓ�)��xѵ����P$��9;���M�nܯ��LD	̻PvH������v�M����+_Wt�����Z��uA]�8�e@�΁H�I13�NyK�/_�/֎���1���]��x�.�9Hi8�7[.�2W��L�*��L30���J����+Axz�[��O/Z��҄U,o����Lt��o{��:�;ﴘ0���.�lS�w�t��U�������C��N�+�$�2�8���~�GTKkn���`m���i���Oˁ��4%�v�L���a��gC�k��:�����a���"�[�fm ��2:�^І��e���*���xuy��8�ɱr6�zWJ�k�4�(͡�ѷl-`����^\�(�1	6�ǼI9L'0���F��(�(���u@ �`g`k9��:ځ��2�o�'����i��'�iw��<c7�X��ᡤ���B����v�2L(#u�ܥ�yRP�_��׻w����@�X�w@D�d�"���c��-���zf�.�Q�!`�0mmFɇF×���`�|� �r�5u`x�_���Ӄ�/;�хD�w��I�t�C:��$�Րe�����0�o|���oۭ��#�<�m�������W�%=�]����/�hMq����e�^W�YF�B&(����g�K{srft�wq :|�_v��0Ϻ���I]C�V�4�feMT@z���b�9IK2��!-s��1O��_KU ݤ?yr�-���֭m]�(��\L_#��"�m�&����m�$8���Г��`T�^OkK����58iu����~ͣ���c����������e���Vq]=*�6l�v�H�!�ͪߺ�w�M��_|��cO���k˶��d}]��5��LU^_f�ц�n�޽��%RO P%4V㋬Ci�Kj�� 54�����a
��1��S��l�*�6f�洬��L�'fge�^�*��,�<��z�0F�'��9�5*`h����|���Ql���5;%Q*!
:H�TX�LlѰqn�� �U5\�����ƥlɶٺu��2M��>1\�R�r�9�)�y����²�1�k�%B�q?��fm��6�@�J_� ��
��0"�� HPV���f�}W��N̆e�������=W����}����c���|��Ev�)�����6G+,�J6���# Ȱ�v2+�N*bjp)�*�C��,B��X��PL�:�͖�����W�̕��c4��( ��������5�pN� ����/K	U߼�^H�//�~����c�Y��r����T�x�ZN��IQķ�[ZE-,��8�l��Ҁ�4��V�Rf4 ��9�@�'�9�H�id��!b�M�xi�#W�800�Fi���RNz�2���]��Jc�Ų*X{R?k��J{�wI�!=���d��3e�.��:�-�f����z��nld�:i��В�� �,�Æ��A�l9����L0*{0 |؜^�e����@E&FG���� x��0b	Jv��0|cv�  @ IDAT4
+Av"u���̀1���*��!��1X�!n�Ӵ�����C��:� $@ۿa#Z�nm�0��Q ,��LN����t�ca���wS㈼�o�襤�c:,��=$���e�ۼ��tߠc�H2����K2ϵq�_�`L��%�!�N[�QG���C��6m����C�P�����f
�~�a�T�HUC�onn��f�H�h����x���q�A��T7p���3&I���~�fķW���LbN��^��9q�8�a���A��`���K�����9�2eh:��~�/Z�� x��w��Q�ko����������Wn�g��0_AK�C���>c�2�]�ҷL|��	�]�83��$�6:�����dO�f	��,|2�X�Ӻ;r��yoL�G��J$��j�N4�Է�o|�>���G���Gݛ��˨	h���Arjn�duL����%	0��%K'�)`� �V�w�{�������y!déd�E���u�����?��>�������{k2=�4a���S�ҝ�h���MQ@�#��s�e�������l"����2A�+i���bb"35 �l��׶��!\0;;�qw����e Q9	Ti\Eb�09e:�$�(���c���@GZìY��h\%l�����=V�9��ɛ��2�m�	�S)*><�T���E��X��-]�̳w&�K�j����~�=�q�\ŕӅW�qk�������'��ɦ�q���7e���ӆ%�3և6wA�RC_�Dt�Dh?67�.��;;;��1��6k��� ?)BTKIb�ō��������Hq�/���<������?�?�a�#u���'�X��Q�E?�M�h= FP�I���a��W�K7j�`	O~��v�����<���
�uP4�����Y�wE��v�ʛ?��2�Ǣ��%L��_v������|��4�b[V�*�z��OɎ*>�n�P��7�s K���ҧ��lUP��j��2���V>P���A�d��Dm5��mp�(��k@�'HY������,'�{���J�r�- ��Q;H8�C��,?jB�B�?�J�G�<��J��b�J&���#[�M���JZ*�������s�>�9_FE�I� m�qSM�0pX��2�C�ٮ�"�5�"�ͭ�84�M�Xsr��6�jm�`�a��-�hOVo�`k�j�,U31b�![p�!ǖ� ��X$�.��n��et�hR;!�&���� Z���zB��84����L�S�����b��L�Sf�檈��!���0��TǮs(�`��X3�,V��aW�| I�Fj����"[�?�R}t�� ��e���6�Yŕ�I�A�a͗ ����py�9f�x#�NY��%.�,�D���^ѕ�6 _RG��� �w�`Y��ihm�AW� ]�x	�~vn�a��:�O_���L��D*�$�x ��gLp4�c�x��z��f,�����-+&�9�9)#�4l`��FL�6:�he0�2y������w��S4	�s"-�`�H$��#`�dcݺ��Ҝ����0z�������\�q��:�^���r��ૄGg�:���"R,�7�(�,���:�����on ��߹뻮@��=��w�vH�gΌ�^Ƙ�7	��H0��`�A��Ė@��Ib�J���`�p~�b�������Tˀ3����6�4W�����rd4X���1^6���ϋl�҉�h; �x�f!���ֻq���Fq�D��Bʚ�l�tA��@����16�K�#\D�
Ȟ �I�]Pw�7>4���(+M��#G01ã��oؐRW~�'�G��o�k[��ѕ���U��'Ən6L���ߊ���G��g��\q�L��|)�.\�V/-&1~!ʩ�[<I�6��E�\�c#�	9�y�/�b��$�h�-_�1��/������۬?y�6y-i����j$���?�?/�~�-}��,��-\� �,
?Z"��!����?��%���-��/?���G}c5�T��LZ4�̡P� d��Ӄ)��l��G�*�!��X�G�����>|�
v"[C�V�$R��� >ɉ�
i3�ˇ$�.��:�Ζ�T�y8/�,U9�9V�,W@��0m����9 ��T�0�'�y�\^]��2a����#��]�='��8�X�@�1z���-Rd�9n���f��#�$~U�P���&XB�l2��.�y�H��#��q4`5��31���I�C�V�'RN���MP�4Ǐ�	l�4QĢE�еg�ϧ����,�>z ?��&�-TVQ�"cx9�ܖM�&������*:eFWկu� ��s-�bB���4�T^��YVe��)8���y�8�{�H���,;�QI3�v0�@T�$f��y)΂e��lxc4f��;y�Ӆc���2�|�U4�d���A���}c�����Z�]3���#��:���[vlw6���¯�$�|`d�)�\&[r����⅍��2�"��r;�O7[oK �4�S�_�C��9hZ���1b`�5"(��E!��)B+��YV�O�$�ǣL�%l����ON�#�F�!�D�{k�m��}��Q�����"��3��	�� \Y��(�0�<��vlߕ줠��C� ��>{p?X�z�Ieu�Gw�f��De����N�J�aݐ:�N$7�R% P[W� �j} MLl�W�&	�]��GJ���P#��y�ڪ
�P0��XW��1	B� �Sy]]]��H�J���ż�裏
xi��4�oI}�����c�j��������3pF�.Ҭ�u2'MU%���s����q̝>��f~��F<�k#i��c~���4�w%+�φ�)~6\�?ɓM�}W��2��
��ł
�9�S�Z���NY��`a��.W<;�BG�FM6Z�1?>l�3n��1^���cX��ȍ~ѵ0��=+^&}��e�Ű�_a�s�)Na��x�;�;;_��\�Y���8rc����4?���k�͗81�a�U<+K�J K�#^����E�r�>_�E�~���*L�c'�8�u)�J'	S�GSP��yP_%/��˟��ڮ������g��Bj�Ltj{�ڰ&(���z
s��PW[F֯�F���n�d[=�9�uYŚï	��������#=:j�z!_~�)�*��u�E֘�1$01�nm�ː���[.#�m"�0k ��B�Q��Ҙ�)��Q���jp5`g���
�Z�4l�r� ���GL��Ľ-�f�i�0pU�5x�; Z�9	�c�qU�B�I�p��T�_��3����>@IX\����F@X�hTE����1�Q�AѪ�?pz8A/��T�_!�m-:���W6�D^[@�4ʚ�4/�161J�"��
jI����/e���-��|k`<C�����Z<|bs�:	@�R6��?��CI�ANp�T��d1���
�P�d���ɔƞ�� �6�))��t�ٸ���k_����m���%_��?�O��ɧ��E� �Yױ&�%21Z�`�"!8e��x�~��k$Y��\l ��d+�q(-��ƌ�D��<ZX��F�#?!�̏�+���S�_bq�I=6dtS�@ꡃ]kk��ڊ�54�5�B��?�	ȧu0�W%91�3vW��en��^����7�HX��Lk5�� /B%33�~��@r�ͻ��c����}�1x���^M~�w]���Ew��L��Ξ%�~�Cott��M}��Ւ�nl�[:�,|t�\� R��$�t,��P�d'�1�{޲�h�k��_�׹+��f�2��'IN��pW���	L��!aؐ�2O��fӘ̓�y��/6oQ�Df<~���Km����f|m��k�?r�9�6�pPX +?���Z��-%k�,�{m޹ŝ��>;U�Q��y��ah��H�E�J�1q�w�.a�$����k�c>Y7�g|Ϧɾ��*�V�(��OS�vQ_��@��V�t*�mmʚ�0�iIYǧ��QJ�M�P{R'|��ˉT�tc�l���|�
�<1��%�������6��>��y�r�ce�A�9&��	`GFگ�=߾lʳ�1�m�M}��&��C=�iX��Eq�Ut<÷%�(ڮ��pH�_R�]�L�V~ꕏ��#��lҸyW�K�O.��k!�ҫ�|�?�/��V�A�L�c9���?�h���,1��C9�#B\����	9�IutȜ��-����6ȗ<ֶ��]��ɹ�P�՞���˾g���4Rqp]�K�K9�;S}������kXϨ3(a݊G����K]�T�`8㩹)WO�a����p�n��4��H%�E������}ymY���'s!��JgL+$1	�,,L�ʥ:ɂ����j��m�KDU(5`���4\��4�<��m��W��҂��|My��'�9�#	�K.���Y2�C�sG�e��|��6:�5v�e�
�V�0!�)������p�s	W��� �C� D�i�"`��I� �P��4d�E|@JI��@"�*�\ɗN�+�9�4�P�!�RHm��p�& �6ЗR�X�u��ܸ͍�q����
�No����U�rP[3lT�����<����]�a�e�r࢙�RN@�X�QO�3�a�pS.������X`�1S����Cjc�)į ��� XiLS�tE��6�w����4
�P�>���w���E�~ׅ; (�t��Z�g��^���d��b�V���&&&��e2k���~����}��I&CNP�r�n��Wޚlڴ	+:��is���w�)�ˮ�bxP�"��P�JP�)�/��wo�Ys&�3"Wq�"	
`��,���Ux`����������ډ�Ic0�g����pIt_ ��,��X���>w��sH�����zߌ��k��ZZ���_�*��A#�K'�֜�j
����tRՄ��b�X����l� �UE�1)8�oS���ҥ+7.���KA$P@������o��<
��җl��d��b�f����+Cq���)_<I� A��A��L�f��%'7R\$�0��q.0�l<4"0�n$?*[�ZaAjM�[�di�(�:.�;g���_|�i���1~tc���?�n� <C���s<1Mp���x^�����~v��q�+,��!;�����&uu��+�+?�))��wMn��n�(�㯍O�+��XgsA��F����&V}Ī���
��N>A7�i
��ih�53��%��G�ż��m��,hV���*u�*�B��R�e�6i��:����JΟ�S��6$z8S�"G�� �Ǎ �(��U��-�l�X:�C鵡�#)S���:~$599kR�B߃`;�l�ψ��!C#R;�l����ؙQ~��@��-d�rb�Th��x;�M��E��v^e����'hl��*2�C^D"�l�>�t�X=�-���� ��j�z���@zq� 7a�blbƍ@bC��q��K��J���d߱D��X��lt�2��m0 *򳋢�D�ɠ���h�S7�I����-�1��bC�́�q��`k�m���b�LB!1���pHv����h����$TC�!\ꁴ47���i�0�Bb��=����;q������7����J�܉>���Bn���d��嬴���P Jy�H_��%�&�O�H4.��Pb�UM��Kz[[�����ߎ�[^y�8r�b��I����Z������FXkx�y�%�uG��$y��N��2	 0?v��'	7I�O����!���t�GO<�>t��&К]Wa�����IU%�J������%y`ǆL�LXh��܁��C��!Â�$����)444t�I��M܀�`k*ը��U՛����߷�=���T��tN���g�g�g���٧������}�7�=�(��@�I���� ���-5�hF�$�8�ĵchS����p�����ŝw,����ſ(>��3�l������kP�~k:��<��T�T�f�OUܿ���:UvJN��u9ƪ�,=�VlǴ"k"�d:�$�8G㈋��e����w=�xVr�Lڢ���:FJyB���;��������o6ʷ���P��>uS�>k�3gNq����<Dp*u���ycc�'6˷���'�B\ׅM��|�����d�>�=}��4&R��uD�\	E���h={�X�H_:����n�h�Y�\�5čx���#~��ӛ&��a�g3~3��&�ٞ&��$�)�nvQ0~NLL<���d�Đ�o��E�r)_([bG���a�Ŧ�`3 ~����]���_�)���ٯ������A�"h�����5�}�ל�q��K�[.\�s�iv6W�6��1��$�C=�B5���������k;�7s�-��T�_�1 ���Q�ft��;��Kɬ`NP��e�l���*�����+
+���H�e���&�+ ��+@T隿�p%�R�w	� aܐ������}N'����l�1�9.O���G5�z���up�D��?� Q r����'`��RѰ�B'��ع@FZ7I"�LI谠֑�3et
q�5��QTŮ��0����s� c�J�(|������yy�Þ�Z�D$Ǣ���5�q�e'��ĕ�{#�JCI|��Wrn��e�rҬ��x6y�{����̓_(is�C���M�v��"�t�ԩr���PPݿ�h9�xj��4�	.w�Wg+�'�E�J@�Hވ��'	;�M�8��*��� ���֏�&�4B����p���-hE����8�F�r�$&-��y���6a�p�ڋ��4����s�Fٺ���ˁ��V��tdD�%#��l&tO�x����
�F��á�PR.��i��t���S�G��+ʃ~
�:��6ڀ�G8�Q�V���D��TE�tA�㏘ѕ�1��4X\�5GӉ�}m})����cz��|��}���;�@�u"S��+�|�m_������g~�����=���Yۄ�����8<���<��Z��e�Sy�Mo*�G��ML<��Ӵ
删?��3����_g�.0�!���!�m!�]�"���$ɥ���N��,���	�TM�<n�����NL�Ty���͘�F�yk�I�m�;�4��|�� ������o�Pz��c�!����g\�s����KvG�{�;��|���b���ɵ,�/�w=���?��w��Y�Չr����_����x`��\_zz������S�jݘ �F����g������9�ÿԳ	˸���V�a�����&�g5}�t��CY�<�F&�~L&:��Xx�\��6����3nv���_����3����3��|	�O��]3����޸����g3M����ir���e���`W�
�ֹ�[|n�ޏ�Ϳ*����EV~�=�iU��̟0py�ǯoUl�V5��띟�@1~Na�����l��E�W���D���p�Fj��d�K��ζ�ǟ�@�Z7�2�? BJ�X��r�3�p*Kk����2���@Qo�yB=9U:���N�@�TǸ�c5���u	�n7�hN%b�m���w�eO���J����ΰ��*F{wǮ�)��qy��(F,���"���H��x*N�����:����m���{3� m�NQMB&RY��/"�"VS뚢R+��`��E�5���MePe�] f�_!�Ұ�*'��{V�5�0��r����lc��bo#��zCOK���!ž���K���A]�b�x�Ʈ�{��>S$�E�\���=w��eϐ�觊�B%�Y�crCHRo�,�4'5��㉑N�����0UZK��6�|�/�%��pDG]53�}F�qo�b��&�U��J�"�k��8�����U��:�Ԛ[�9�D+tr��3ZG�8��e.]�F1u�*'���={w`�q�b�:���Pt���<V�?��ǟ|�+TڈW!8�n����hf��B8G��+)d��C�&	iIQU�&�yN�����X�� �F�B�^X��_���g~�ߡ�4���i���)��/��8���Xr�O��%	F��<�M4�E�<q��x����8���W���z��O~:������9�����cQ#�aynK�q��@���r��D������͜ia5����zk:#�2@ο1�(�o���ŕZ��Z�g�Уb�B�j\uմ��0/�wD���f �_h�o��o���������w���k�ݾ瞻�@2�5���iE�Z!nS�7�b�ԍ���#h#�����.0f)&�@�t�*��p'7�&\:Ĺ���ku?�ps�����_�v��UD۫S�/C�m�����3#���v��׵k�t˄Aw�Q�e�b�M���	6�SDوb؄�v(dC2������0�Y�����X��y:;��a4���ǀg�v�H	+k���f�m��Np��F�E���Y�\x+�s�����g��4z4�;/��q��9J��?�����<Ԃ��󯚮фU����f���|ϵ���W��V�8(�}h�1g3b9�����X�י�6�\f��>1��+�غ-��Z:T��&���80m�R 	�꧙g p����H�j��@��{���H$	X���,�B?�� X����:�`YR�X5�KU:���K���A� �����
�r-*TȄ�CO�k��<5��:�lU��@Q%7��x��g(���*R@�v�����(�*N� j��/�boV�k��V|��E��@�\�rq�mbfԔ��4l����E��P�8`�,�Dèm�0�.iX�b9�1�n��Z\�I&+0
��[N�^���ݟV�P�{�-%9+�;���w�"�m�P�9�L�������!<�H�G���V�D��9�F�k�NW�H&�����!"8EFk�&p਽���BS�~�=D����s��d�GW��ǹ9v޺r�:��#-{��@8v� �X_��F�8��Q�b	N�'o��r��;���8R$k��߹����A�r�E9��v����6�.�m�z��f,(Z�`���i`-(w5r;���MP��p��� ���{�FN2���u_���P=a=�����-�=Zx�].�;�
Hb���D2���T��K�`�ٞ�\����bX�>��i61
���W<t��?}�ӛ}Sz��c�`���")z;.�E�=N�,17-h�� `�^��/����r`[�~S�L&p]�b<���21���b5�?^�@��W?�^��$����ƊnyQ�.����e�&&��dF�:S-Eu'O�h���3�[�p�� s"=8C����p�*���ލN�<��%��*��N ��D�� ���ʛKKXz�<4:8ph�k��49-����nN��2ĺE/z��֦�M��`�@��N�l���<�m�w��A�RH���h��@�Z�}$��a3����S��&�3�I�X��ԃ�o�6�9M$���c��Z�ݖ F���� ָ�q�"aʚxk�����3C�����tԑ��ƚ��
�j1�{"���%�L�Iv���Yuuc�i��aY<���ɉ��v�%�[%�U��2�E��D��GH�@�իx綮=����k%6m��̜���ן։v���VG���ȟ�2�:&v`�ٻ�Ϛ��I_��Ѱ��#
�R#*j%���;I\46ӦD�8�nP= �³�Ҩ���m�Jo"GYy5��k嚟���d\��
7@�Vu�c{�C �d���[���l̨g5�7����6�ك��\�G�V��O�xq��F����h��G4ꙣǸ N� �QO�� !L���Ovx�H��Y��b�f�
+? �٨���P������M�`��[E�8��c��M�db`y@xV	x@�#>HX�<�X�m�Epԏe`��*R[����FM{c�,�?:3�\� "b�Q�_�P 6}N��P7�*EW��
i�G�o��V��]� J��ʼY��ʶ.Zޗ�QhD˅��P�`Ƃ@��t=��\űv���JX�xr�ǅ�}z~�ז�ZC�,<YGyQ(�\c��-t@�mQ�B��s������e?z� G������.ɯ����DV<�UO������V���vF�V�_wgNw!���]��8��Ǳ-�8���\ت�Q�Oy�<al)�~�nW&T$j�P� aםa�y��b�����%8K�����TNG
�	�!q�7��KD�]]����^�3��a�����l+]��V�A�����6��
��%C�s�rJ���K܆��us���~9�}u���q<B������7���46,Ҥ��yG��n���µ��x%���I�@�d�KZ�H�{�5�i�]���ӧ�?�N=#�^m��:���.wN�J���g�]�i����5ק�q�����BdF���&!�/��^x:,n{Z��{�Nq��U������p��7~K9��o��s�ݳ�ؽ�8�\��b�(�&ʿ�>i���70]ibUT�!(ڜ���]�x��52O�mb��{ݰ��<��0Pɵ*��E�����ipw9��)]�t>uKL�� ��`�X��W@�	+�b��c���^8��Xg^bw���L�st ��r�	��71
Ag��Y�B>����W�ʫS�
�FIׯ\.�a6a�#M�v!��`n�t�,6"�&)ӄ��8ߧ�.�䂮A�-��7h;u�$^5ap���ЗR��"yq���4��3jk�kA�,�Ŝ����:�XQ�ۀ�\�X$�M⇢:Ď6�`x-1��uҮ���N�s�=�Zm�S�60���{Eu�K+K}��i�p�p���ߍ�L�UD�|�ԡ���b����p9��q���T���R�is�L�]&�D\O_�G���r9����շ���O(���ZD*�0�D���0��p%|we�JV� +��]{o���ߎ��U��_?Wq���ɑ3���D?$�x �� H'Z~qe�F�{M�#J�<�m�׫G�����m���|n�y��g]��ֿ�Z�Xu��斺���;W=� ���,:i�Y��ߑ?0�qr�����|Gys̭>�[��MQ#�FV-�n[�ʧ���ǝ���^��B����b�l�����ĸ��_Ȓ��6�Q.�u�DpٹWǋ��a�U Ac<��ER����x[�����E�Iw�V0�r�Wm@�~��R+��.]��2�'8+�{����2J�|�N�e;������\�Y��oU��Н��&��Cm@>T�b̔���X��~�1���հ�\v��Hq�w��3�/��av7�,�u���BT8�7��M��L�R4t���KR�]�ou���y���?�~��~6b[�������m4;?���{>*�cx���[]#w�Ь%��c�ǊD�D i�R��Lf��Z�y��<��A�2�z��4��&�<���J#���ꍛ���S\��������Ǌ��P�	6�p"�1Q���KW㾵�+S���%Ƒ�&�Z�d��0�u�]�t��)��������eկ�>���Z�����8�ʙ���;�S/�,�<~?�8��ey:C�gi/��qiYYc��)q���V���Cw��/�Q�q�,W+&�f��/ˢ1I�xG\����mr�h����8p^�Z�؆k+Ǭ$�2@�X����'z�P��=�7����q����x(��������MM���Q��/B��a��X�0=��?�\���*^z��)��5�{q�:�2qd�rl�C/}��~mz��B'L�ºxo�ɓ'ˣG��<p�Ҿ}�gp�.�*0�{�/ݟ������wa	��(�������+	-�#�9�|P�(!f?�'����Ŧ��s\Udy���e���՘=!~�N��G2�$��3�����or����B)0<�]���k���c��"��sOE��ah�Ť������c��"˸a!4�w��߅��^G�P���g'����$��G�N�ʧ��d'�mq�lƏ`;�6�O�K��;: !�&3l��i�H��&o�2���;�����9,�m~�89�����m��0���=�� '�8����s������+è���-�N<<�=�$�߈�2UQ|U,$�Vݞ�U���C6�Wg�װ�2�Gj��2Zv�3�"~4D5D�\1����{�#�$ry���&"�e�&t��C�x�D�6�BO
葈�zk6(�V���<��J�ᳪ�#VO���0R'D"FQ�ʱ�#2z-���8�/�#�e����at��/,�A�aOF�
�4��ԍ@���$ҬgW�j��ܩJ���e^��'��r���F��S�l��'�ͮ� M��-V�Y_�����Q�e��	��D�P���	B)H"f=F��_F�$���S�%�
_�"����,+��[5
,�obb�kI&rS�?�'y�>�� y��,��ק���բ��pY�D����K��A�bc����All��q ��o��/d�t��rE4Ll�j��{V+�O�ƽ�|q�@��1�ACı�.���Ъ�:s�b����kdO���D_'.�p�����bd��;���&'F����7¨B����c��5���Mӿ�D���`z��G����'�Ҿ;��9��Y���CǊCG�P�!A,�K�ž��K����k�ŝwܑ�8%9��&�X�Z$D�X��9���fl>pA���s�����\\EhrQh�8ؠ�0ǎ1��$���vƿ'Ӣ?�'@;Q����M��;���B�C�7�\�|	��\��t�����,F#������By���b����'��� ʂ�A����u)ʏ-)s�1��Y�c��p�!H,�}���z:7%�]z����~�I�XO�5�����8q"r��)�7��M��c2/�Sa�*�>}:����d���(���&�����<�G^�A�,��uS�.�Iމ��K���V oJ(�i�V�L��s��#�A�ݵҦ�S�p�a���$60��펍I	e��m��Օ���G�z�3�?�$��*F�|�oJ�"�`IT#��x�.�M>�p��ʷ�#�AQ��J�F[U���6����prX�f��I�ﶛMDգ�sB�4�}��fn~7���!Y[
�9���4F�/��߯ɣ��¶���c{:#��r���=n|ۄD�׉����o:F<�я9�Vt�׮��WLZg��~�o«���$����0y���32�"�3��"D"D�)Q	���b��%����+ Q_��A�����GƳ�8��E"��,r4���?H3��e�1v�Km�DT�� +o�7�]_�`W�3a�?���OK�~[GlR� ����²T��s7i�V���~q�
���Ƚf�"d^����Q���m�(�D}�_]w������jց"����"pS�t�A���D�U��6����� A}Z�Xݽ�7�i:�V 0�h$�h)�KXӌAb���كy�h�Ac����v���ŸCD�
�9q3��ol��1�i?�v� hd(E��&d���)����*��n�q���Nv����9�"��y��j�.s%���b��x_:�qO��86��\�6ϝz�(�����V9���� �J#���˟���VN�=�aN�M@h� ��p`�j��z�3���te�z�xq����9�LWnpu��܉�
��qB��2W���c��a���hJ����^lîAXpJц���<*��2��nVQt��[��wpu>�Ϥ3g�qμ
�?M_8?��s�9��� ���#�a|�Å��b�i|�!Ǿ��R>zWq��+q�Pn�"��ř�ꥋ*�a�bz~��1��U_��O�'�|������=O�.q�сC��N����CB�9��o��e
.��\���5	�6�LK�D���[�7Q+o~��:m^�e{�'�w�I��Pz�Ǣ��W�g�uԀu��dY�������e�Xk�n-�W�[?��h�cd�j"A��ĞbA�2O����	�@An�	��V��d�	��IݸCX`�MÊ�Z�ث0� 2���ckG�@�515�>1ȯ"n����g5{cg/�5<s���=��HB�����2!{�!�d{!��[�X=s�&��{�� ��V~�|�x��7?�5xZ	]�b9�iU� 0�Н�Ux�Kr���U�Ny�"G\�#�8U5n��a6a4ߛ�s�엿����>o�N�����>b�4�p�޾�JF��6���o�mۿ��������&v�B�nێN��Vws�)�,$�_�4�V�j/��2���
gξ�1/����OV�.NUրT'3��uD��}��� ���Pj���Q1"gǲ�����v��ѿ�b�9i�:�#��y�G&x$t_ ����x	{�0�5�e�X`�#�
��!��pAԩ��{^��S�"��/,Wb58_�T�nd"	9O�`QK��<gK���_ye���Sq�}�2�
2:"X+���[�m\���d~���C�>� #�T�u&j���˦�Pc :JyY�Pui�q$y���'�3�{~K�V�똮ƾ%��b�A��]�Ù1o�
Y�E�"^_dQV?��h�
.�e�."��:��e(�W��ے�2:Mދ����l]$������ЃG blF�b5���S�MN�\��*F�{�N�&foRv �wТ���:{Tp�ʮӒ37Yk��]�J�X�U����짊���V�*���W���X�QP���xO�R3�r�i��J�4��c���t�-�cK�Pz���;�.v�Hׯ]ƞ�2��P������v �F���}���%�!q<2�b�@|��ٌ�����I�� ��p�%�p���6A�������	!\\Bk\�b���F��<��C,��H�8��J�4�����B�ַ~e����qJm�D�U�@���kQ�G|���U�l��U`\�x�A��=ww��h(�3���{&�7b!;J�׶����\�`��$T�s��Ǻ:B~K�m�	/$\h�n�:-�A�!.�TB�ȕ�����G>��v�)��p��?�����Y��(c����/�2�I0�گ�Z��<8q6x�t^�!�<��B�%�5�()���r��7:�G��>��o�C�	��N���IYYt\w(c�O܄�-/��
�l@�[�](�ͅb'&��Kr^0K���,vRa�0�%@[!��a3R=~x���_��>[O� ��%��IsV��7�"�yR��u^��%��u�kb8���H������7aW���BT��W�� ;
�|�6���׸(������u��L�|���/ ���m�(���T��>�E?D��f�G���:u�;�k��?~�N���"ë��3�6޶�|ow[�/���	����T��&��a��G�'xʽU���0��E��H�-~�� 9���WZG��R�
l��:�<<h:3
$__�Q�Y&���<��]H3?�b���S���(�1����DRO"9�\�����厁<C7�}��Y+�@1i G�:]�_3pwO�A� �>�1d�o�{��bݖ��*�(V�C\p}z��^�1���I�P�V��*_Ws���r4�f�0��H����'���V1~)Vh HA�\����𔟢�/	#��L���	��bf�J0���-��(.pۻקH�{2K��e� 8&�5ǰ�;�.�x�)a[Hq�F�W�@Ae�y�K@�����kAi��Ģ9�3r�l.q)2����ZZk��2����.-z"��Z�˘|�Z�#�?�mW1=����wAŜ{��0Ű�t�T���2sJ�L������6>|b��O��Nח��ee�5��P�Rݢ�nON����3s�����\y��E���,w�$9�)G�5��;�	��5B[����}�����]nR����7����R�<Ư�9���;s�fD���-���~��R�_/fne+�q���>[<��3�7�.���]=�;����ر;��Y�A�O��=�ɽ�Z'O��1����p +���QNɱ��D
�Ӂ~꺾t�ks�<'%_`�\��̆Ik�]a�y�7����3�) ^V(�4�7e���A�.�
����K  @ IDATZ��á��Y����nD����0�x��ѣm�*���y�����jל%9E�r�0��T0\��õ� �  @߿,�;���`�"w1V�Q/�K��9�1/���&#��b�
Jck�M�X��ޘ �L(g�N�����&�@��Y�$\>��Մ!�v�	�FUh�Q���U!������1q�cP�	�I+�2�<�Nd��ƣ�d��\�i}��~���i����O��s!�ʨ`E���,X��me�p`:ޫf���������֌S���­�Kֿ=�m��~����<��+�N=̰x�� �zk�����g���#�W�0��"r�f�1@wV^��Y��4`�i�qM8t�~�2G����&"An_[��/��fUT/�ƻ�x���@� � 	�Z?��7X�V FD���Ʈ�e��*W��|D:�s�>�\�PGp��`��F�E \0�����N����,���QQzkڳ�F+� z8����jD��AR��ڔ���J��#u���F�-�������`�u��� h$�4����-D<������x������V�S;8^���xj�G��QLχ8ϸ�r����� ����X��G3�On=oKEB�N	V0�M���؝җ����h�6"rt}�����q�� �+���\P��IXp�#[�7J =cO�V,��6ז[�r�P��$�\�H�)<�t��AάA�R1�c��6���aU��T+p- ��T%�3cܗ����A��J�鳮�PC�]��2��GQ�)�P����.V*�I�����z\��=�42H�Q�����U�?�Q�#!��Kʝ,2GČ8���G�,ޑ��8͉8.��f���}�+H�m�q���b7V��������Ci�ƁhAN�q�{��@�2}%��S��EĎmD֫E�����/��EGa�����/��l��W����(�}����$����2
Zq����BQ���X�9ʩ���ph!�� �I��ha���i|�d��1�b�[ �QLgN�K�p�@�@���\0=��n����o��}ߘ>�}?P8���ЍHuQ!}C��;'���W^J_���\�;��W��bq����p����� �1|]5�DVх�@)��Us&�7�8�H��4�.rt�YFg�aP7�K����=ۤ����Q�D{��#�[dKhM�"i���f41��1����W��.��I��{����W._����۷��~eW���pD\q�����S7��E��"��*�D�?e���:jR�ݠ�@�bG�Ǻ.�i�Beg`��i�jQ��~�iD����l?i}��*�.~� ��t�?�sx~V�L{CGf�I"�)�
��TF�g	Ef�W�ɷ�5�UiDNuB�L���£�nx|�jӘ�Z�"_	� ��lP�#%��N�,~7]3��q�w~���`�]3^�=��g�݌�.��~�x~��k�k�o��ao�i�4��k%�n��ɶo8>�Q���F�GxFUb�z���,�*�-?��5_ouvw�u�YKP�ÃB�D�����X~p�DI�tY A
��G�!��ݘ���+��}v{����Ȟ^߈���]�����	S��4"�k3� 3J��x��T"w〔LK��e�mz�$�\dlO�`��bE��������eN���Z�"bw���n�\*	@I�.8B3h�9"
�8"��(r��$�q�I�k�mH_�9����(nG�[F�!��']�5�⽞��}��O)����'����d��#���Zt������K��X��u�C$�p����<���'$^q�c�W7hAX�h[HÈEo�Y������k��ݜzIg��-!�R�ztr����^v$z�	�P��QE��b)4���Q+�Z���F���R?0�߽?�L]�r+3�������O��C������g�C�<�ɲu�6��yt��9-6�©��j�@ �.m�l��;���(EW\x���ΕK�FIӉ���2�@u��\alm�Y�*��?{��rn�<r>TP��,McDqek�69���=��~�-HR����P�m��j\c���b{�dMy�:�<`s���훺z5mb�{�wA�$�Ư�w���ԉSYld���V�H��q|�;���0��z�x�����p��R�߅���V�+i_�/N�uu��ɝ���鹴��ݩ���=Ŝ�r��u�!��,c�4��T�gz�G��{���U�`\�Z��~�<Z�ȏ�k� �ou�8�;����7E����3��x�'�a��CT�1�{����Iu�����\���2�Fġ�X\��8"2[ �h��4�/����	n_�!S�K��Rr ��粰K�!%�KG7�H�b�k�v""���Pr!]t�iZ�X���F�'�ĉH�g��~Pv�����@�˲s@뼞��t^ x$ˬO���&v|�}���:����VGz�V\��(g,H�ޒ6"��uQ-��w�+�-��l�h����($.o�O��� Ov�>X�;p�R���������؊ (ˏ ��������_7���,�i�t�ׁ����lv"�KU0~�=u픯�GM���"�"��mNs���hDh�m<�����[4�M�z�0�%"t�b����*8�l� ]Q�����p���(���<�E�L�5�d#<���/�X7�Ё`���G�*�^��Nss9��s[� ��^�q��T	CE<$�2�f]!O�����$Ē�E��	�
��b'"7	7�o�+�i���ǂ ���J!Ŭ�c�t1b�PTA\*�ɕ�Y�RC��E�{�2G�Ӄn��4�]7��O�у%
�*����G�G{�|��ĉ�����#ǺqѾ�C%��+p�)rVG�D=�`��6P�fE�~Z����N��/1��5!�S(܊�CF".ZC�|)ч���gKKA�3�+���e�.C�Mo|��k�ŗ� ���ǿ"n�?w�Rz�ŗ�4~r�$:wc�av"��Զ��I����q���hǉ�G�Ҿ#;R��$,cΠ�v����b}ᦜNK.����D�ć�:/��׆�YÂ��)˵�b��Mꆽ���X_+F�����b��]�}� "QZ�i������9tl�v���K\�g���B�����k�x���-?�CV�:m�dM��^�r!t[�48� �����*P�?r�W�Lp�����+��7�?R��U��o�f�����F�Ǎkj&��V����`9u�b�?�'��y�/ryq����n�?���H��n�p���fl��}�Ð� %�$�B�7c/�߹B�8��s�	q����bnu�\>�~n.C�����Ka	�R�aH�i�s�y�h�J}۷}[������,����J��9��щ�Sk��ޘb'��-d~�qi��=NXL'L��`2S�:��t�h¨�r��۹��v�������=������S���h��i�����o�u��e��ڵ`�@ /j�$V��U��)�_�Fr�4�;𱮸��Bo�b�`�4���}�vw�ac������ڸ��$� ;�����p�ժ�� $oJ��t,76@�ػ��������N����S�Z]]��g���{��fB޿�xǎF<�� ��l���T\�-�h�/�?�'$��|�,�D��A��P_^���LS'}M;�8>��3����d�U��6�i����x��ͬ�g��3��Խ���rE�h���������@?2���&�*8·��i�(��Gψ'�"N ]�o�Z	&vJ"Y6��R��v��Ҁx��Al��8���ml+�IHZ�/A`	�8pB,gALk9Ϻ���S� 6�Y������y
�v�(��
����.�E���T���w���S{�Ó,��K��Q����+E����1����|y�̙�7>G���N��{�@Ֆ���/�����W��<�!��G6��l�X%٧�s�ŎqO�-����G"��0r1=2�qC	Kt��_�a�yA)UI}��	'�P��n"2z�O����?U���7`1y%qEI:z�>�\)=��W����/���я�w�({K��\�1u�]
II�^��`���9��B�61lx���[\*��e�O}�oi|�X�8;w�|�����>�y� � �=�� v��T���!�`o���U���� ۃ�y�/{�s��s�,�+N���P�'�xC����rv�h���P��h��bм��Oiu����n��H��c���
�=&v� ��\h�sWw:sn
�݉bv�M5jW��fyp������KKd؃"��� ��Dm��f��E�om����p���ӏ�����49>������3�2����`$�����,��/�������ѣG=���Qq�=��u�2֪C�z�_�i��8�s^�G� ���6��Ob�����w�����s�����bpdؾ,���.��(M�#�32���v�S�2�B�o�hE3���]^���u�1��ᜳ������3��߷���|/���9m����|�q�f{���J�eLʊ��%mh�8�+�����M�_M�e�\��|���N�#�ƿ��J��
l�V	Nv�<����"jU_-��r�k��lbwP���6^��FC��;n�L��TH0(�@��Ŏ��K@�me�^��R�b֭��U9n�c����V��^��q�U��V^W�
���$Uxn#�}#f��G̿����Z�?���N����G��"m��oӯ�ެ���o+^ym����e��1��*�^�Së&���o-�Yp��8LF�'�lR:��F����6�Pع�L��-��S�E�5���i^�ӄ�;.�^��F xKU�u��� @����"2� ҍ�6��q��d!�Ltʑ��5	)E }�m��Q�^����z#L"��q!n8A���(]�IC:		e�)�/ ��E��Ƌc��)�+l	5Y�}\a��+�+��b�b�,9F��UL�,�����|K�yq���Pqh�]�4��ׅȎM����#�4A���;ɒ�Ά��������X��Ĝ=�=���<W!*���W��3�����q36�I;D�/���G����b�7��J}�uy�d�P�E�d�p��H�[u��I�e�}��������}w�_�*����փ�ki~�k&'("z_p]fQF�,���c��+�I�4гQ\�t���k���=;:�2|o�o�]������g��	�U��s]Ek���G��9}���#=��Ujl{��V�F�w|����/��~���_�&���&��θ�A���١���m1U9<��\�N�l��c��!�=��1%�F�<�Zi�{��<����7#܍���}���[�}u��`�|y�x���r�����9�2�����O�n�}5��������C9=;�c�4F4��0�T��i��'�C�Uf�q��JO��	&�b�O[�7��=�2K��p��"�����W������oRPl%gJ�m�j�ѣG=Q�~�~�X��|��Uާn\K{�Hk�e��x����O@��bC$Iͳb�}�s++�"�����"��߾G��~L�����o��Û �����0��5���&�����o�:LEJ����8�OD����Ď���Y'����ٌ"�W��o}U&��X5�m������!c���I0�ܩ�%����ׁin<-�ɰ�P�~V��m1�;�[� ��%��Kvf���L��n@�{���F2�	Y���z��FH��oU܎wd�����L�ߛi�_~��w��:�V����U%�T�����D��8��89���G�����Fc��w���o�:ހ�E��wU�&̈^�t��w~o��~�i2�u��~�a��g���e_���n��G'�Mk��]'m��D���89n��W㿎㣙��&�d)�ǳ�~��*�����x6���f��O�H%�A.0�jc?'B�Ř�#�T��f"�!��+D:�tM�1�;I�p�͉Å�3HI��F.���1K=��w3o�C�*x�Z�v����'���nq�MD/�fv�sz����`� 휜d���g�}�ȑ����������?�ߞ8Z�NS
�	��!ND�E��4X���υ�ְRǼ]�P2 d8e��C97�.
����������Y����0�����/�
�XD8��A>�^��s�o�d1
�(�C贽Z����c��c�����Z�.L�}�;��ϧ5�����_x��/<[�Ŧ¨�ڷ㎈I�s�2��3/�I�Q^e��tZhû�:��pP}���sߒ>�������$���������|��[�@����% �-�I0��;wy����:��e��
����'��!����C��ٛ�������D�t%���X�-�f�"ͥ3'_DWio����<���۟|k����h[��k����8R���^���[^�|��������_�v������_!aPA���(����*뷸����o���>�>��i��������/���n�5h&�䑻k&TuJD����w�O�
N$��3�Z�����l����������R$a]:�'E�;w�G�sO�����1�w��*�bz�'�V�G�&�Dz��p,9�Ř@�j+O����>�h�W��uş������C���Y���z� ��b�B��1.\�^MB�s���9��n>�o�w3�9^�����is�#?����o�������̿{M�ة�R�O�Yk��4r�}X߸,��	���%�cz'⸛��+e���rwr�wZ`��o�+]���n&
)��V,�^�o�e0.��=�0�`Bg�`�Bv���xV"��*y9��q�W��Ҩ;�<
ւL��٫"99X�/p��(O�����m����{����S��;_�L6
.��3�u�!���+������!��
��W&�z�԰��+෕���}v�k�K';�Że�.��݉��=G�0��_G�u¨�CA�Z�l�*b�=����Y�-�E�������ԁ"�`�O~"���g�A�<�i<��������È�G�P-0U�w�T�X�v�4�E��K��G+W�%g�!ZB������	�J�H�hAh0��lؠ���z����Np��Q_9>H�ԉ�k"&�i9. �������ؑ{�-�L�"�j����u���4�����6�p��>��S�7��j�_EK��������o+�fҥ+�Yt��;BCq�hF\�뽻�ni��	`�˛a܎SJ�&UY�ZҪ�Ns̱/t�-)p͟��\(��x�|v�Ǟ�g?	N�-Px�b���t��S��;��������rYk����g�IrfGͳ}��/�<��\�O�{�J�-*f��l1�vx������'��������B]�g��Rы�G�^�ʹil-J�pJm)����ow����)@�S�ǚ���q��ϟ����/O�U�뎣�ҵ���Qǒ� ��ƌ`lM��n���X2G)ڶ�AK1�A���*�2ۆ�^NS�.;�N/��Jz����;����wP��G��i�s���̹����M]�Jk^VA=��d�����o���HO1���T\G��s�ǯb��Z���R��th�D�KW���g^,�س�8�oz�O$������b1��S�/]���&�q�cEk��x�������.����gΠ+W�_ƪ8sK(u����%��y�c��4���������0���|&9r�D��c��	r���_�U8X̃%�Hz�i�u���29_��T�d�IXi�����Qs�m����KO�c���b��b ��:l7�8��l0,k�31�%�e9Pz������)��m����ö�x��/�/���	c{���/�Ww�/A6պ,}J�V�&��f���9�hN�������K��((b�IR-�v���x�`�3N���B��L�E1��1�[�Z	��sH�^?�?�aqC_:I�m0�o,�Ͼ�j:���or�H�\	��&b�CTJUT =_�v~o��>'�����Ϧ��A�ӓ%����W�/�i�Y"7ʄ?͖	�N���6=�yt2�l	7�����ĭ�*8�G����'ZN��d��WC�ǖ߭���[Vڨ��֭։S�!��O3h�G����WF�Pu�5�cg+vnN��j>fT؜r����}������3���|����bs�G%7�Gz�=���xV��b�PmI��rH��.�Kr!v�lDW�P��+���o:�H�1q� �!�R'�9��@�0ߜ�y�>��JK��~������X4�8�f=��?c����'?������V{ˏ��<�W�:��d_�9^��,ށE�EX�!�\����Z�m���7��E�!�0���r�i�����@Oٽ�\l��x�B��w>Q��_�P:~�I��X����w�%o�)RR��O���{?��]���c�G�⢛������s��@w�9v8}�w?��^�2��^z�������k,��9��r��
�$g�������a�����;e���>�mÞQ�M�ũWN���!0��&mH�Y<i
&��!
(���b�P�t�c\�e�d#_�{����3��4	��k�7�b����chh,�`��z�b�N������?��p���/���;04y�8w�Z������~�Wʿ���Aq�]�ǭ�/쟦��'ˣw*>�����/������i��	��?�O~>����Ǌ��9�y}���ďcG����o)V��/q�n_���A�V����Ig�M�B���3Oc�n*��ǝl�}!�l5�¼SS�ݘP��ut�փ�$���gz衇�y�ܫa��1gQ�6Ƽ��j��G<��Î�\(9f_Lq��q�<�/�N�>��p�x��ߎi�c���Z����BQ�c�9$gvdr�k\<4���QBqAVI��v��ND�x��3�6����o�w�����g�����&��q�a�����o�6�,��(��*2O�A��*���
� �㛪a2žͮ�NXՇ�K��f�����@�&t�4(S�ǟ+B���%�E�w�+�M����.&^���U-,<*�H�3�)`�}��x���oPʣ�L�u&,���*!�ԐB������k�7�������bow�/?�ޫB�N�Q@��|��Gg;h�ή��v�fX��u��ɿx��X�Kn�~������?u���e��ۯ�?�4gM��h�b��t�n.w�&��U�1�;�2�sZ?�� �i�wt&a�*]�'��@�p����X��&�@z����tq����x#���;�9<��h@�.��%�$r@�4�3�S�6N��< N�7����C�i�� ��o�ب�C�E&v��G��}!8Skx*��\m=���Rl��R(�/sA'� �l�[�x��W�v���t����+�ӱ���0��|}u_xͻ&C����j����L���'v�?��ªn��(o�������J!�)I9�RQ�:s lҮ��z���o��t߁
���/��i7@{X�$2�w��j�]w��?��?P|���@y���pQ��re=���<�F0'���b�K��G�w��G��t�Rq���^D��%2(N_q�,����v�xl�9C�K���{X���2��e��m��L�/b�"y�aQ��t��*�p᠖,�p�8C[�i�X?]�kxb'���zc��ܙ6���q��4���N��y	
���Z����gϖ��+νt���ؑbxρ�;�{��5����Z468�.o*�N�F���;�e�O�����C���"�&���0ҏ���~������~쟧������wm����N��L��?���w���Wf��r
rX=#�r�w-�+���R�U�pʲ�n�Gd&�5���pY?��c��PJl��������Ņ���G�G��������E�V#�����p��-�_l6��Fq�I����b��M�F�JXI$�̎^Rq�S�D��SQ.e�|�Rq�����Ѽ��Yu�ՑѢ/��A�\B���[����`��i�
�/+T;�E~�O���Ͱ��9n����e��K}�4������5�v3�n)M�%�T�Hk��"��ZQX���:�̴���'���*F?���U�[�.�?�}tP�9
e �Xl{�\��Ę�B�L�[\�,Z��x������j��AM�u�?�3 k��Lt�d�v3J�J�V��E'�H����K�����lD���6�i���=򏶊�*��5P5�V�f���~d��;��Y�ܭ�������N���O��{~�Q���u��ER�<�Ӊ����$�%�5�j��s�����k�j�u��ON[�G��K�5����i�_��(q��^ӆJ����+��l�M���f�^r���uu��C������ą�r�������_��[� ��jIx����`�7L������SzI�P�)�HGx�W6�#�Ʒ�.,r����|Ϟ='ޮ]�ᮼ<z� ��F�!�;F����S@��B�/��r{��Bj�q�S�(�?AQ?	�ālj��;n�T��2QlW��3��w���-l�3�.���O�~����H��a�En��"t�αG2}��,0M��x��O��y��ز�`��=(�R�y�I���Y���gj&���@ �y�Di?⢞�L�I�X[� ���Zk�i�B�� Ä
]�Qc���� B��8�am{4AC�Q��P�����V�MX�Vdi�<��2\�^N�� ��F@�9���V�P��K��ôj;]��9r��Yq����/��qV����⑴xa�ص{'���8۽k�ۇ9¿;��x���J�09p�cjӘ=��.O�r�x�7��\�����/����Z�9�Bz+�����حO�ai����P]��_��`���?p��{@�*�g�1�QL����� ��������G8QȜ�F]+n�L�'�xtL��y
��q���ܡ���3Z�ט$�(���.1ׂөn����[�3�AEm��;>��X/w�3J.�-��=�)|�����x��Z/��

��Q�͵�N��ʢF6h��C�Q�Zv�Ԏ��z-��=<�i���x9,�i>s�엿s�&����᷋�V3]~�����SF��'v�c;�K�U��A�h���S��-�����Sx�%==��눮�74_���U`��&eoU����$q �heѭvZ|�n���p�Ï��Cʭex�;��u�?��T����W�����@W�ҏ�E��@�nV����m�8���\� }T����9H�Vb@�\AZ�L$�;@��\*��&�؜�`
ɋc1����Wc`��]삻`�rZ�"����M���-����(�]���rՄկ�}�<-wD�� ��6;�`�Y���OO<
`�:�e��*6��'�F��tq�K�x�n%�ުrѢ��U��*��do�5�F�#B�զ�*C%�G�CQߜ"_�i��F��j���5Ԙ�<� ������S�
��"���u���t] ��(IU�:mlL���ԑ�����mY�(����F�r��K��(L�={vK�C	6�z8�o�c�|"ၑJl �"���������m�AKșeز3V�Ae[�dk	B%�҈=PH�*1���r �o��"�pw��;��G�F1���(�DB����6Nk� "�9{DEk�d&��k����
\��W�-��c��x�S�9���<4��V����d��H!=�a��a��Q��?��-6�V��Z8.���l���ⲏD;F�Q-��8ۧ�:���C����޵� ��_��n�z!}�}(��8��;q�?4�^��,�ju����[����#�8<6[�XG�	��x��5�V �.]�XLs:nx��tsv��v}�ؽcg9�)������T�D�Q�3��P��@�409�tea�hV,�U� fBpt}:�C���}���V��\��'�Z�KCKH��}@dT���8Y\�a���e��}Ş�;��m���t����@p'ی�ޮy�=�:��ӂ���;{��i�s��np�������4�S��[�C���<������+�5��bn��\C>�FE*.޼��=�ط�8�p_1����$�~�\:��s�;��H��W�1R�����Iڪ�Ӂ�J$�����������r�Dk)mBx�Ŷ�oF��	�l,E�L�An;d��A.1~�ӡ���⦇��a�4�J̱�"]�v5.zuP1wuz_[uI�X'�f�4���?Ƨ'Xcu=a��v�Y
�G/��2ze�ӧO��t�x��S�����x[j��Ѯ��
n����ɼ� lA�N����R2���ѿ�I�:/�3&�5���U�V��0�G�fX��aN�n�_�	'�����r>���N#�]�w�R�i�_�4z�R�Cr��خ���}1��򉴁�QH �r�҅�~�r���.!Νoщ�A?g	�	#�|�Q�x�����3�0eqnb�ꁽc�/|�7���������:���0�߭է��c���P�5~v[i����I�Ԉ�P.c�8�)���ޓ�
\�5`E���zC�&�+�Gt�+�]�J?�"M�2�γ�R(��ǲUo|�~8���S���7�r��4Lg���KuK'D�\�f��5��.Îv^�O'��忕�����������w�������e�s��M�O���C1��j�N�L	�:7��2�÷!�"q���o����	�y�_�F�S��tZ_:�∻��~7� ������T��uU:��������N񐢊�p��N�\��<�$܎����lQm��*�AT�����	��ȢDYq�z>�MРn����t�2����-��S~�]����U1 'iq@��ʁ�ĸ���<��Pz�Cߍ����vq���u:�>�>�I[_[Lg.\M����^f��*9��u6YT.]������U,�Nǭ�sׯb$qL%�t���(���Up�����8\v7�s=�ٶ��X�������}��W�CE�Ї�/�_��M�s�g�nN�o"@�8��/��\F���s�nt�n��I��#���u1ݼ~���;��-�}W��F��α�F���":������#^�!�J��,����($�k_�mHʔ���[�[��M���n���	Z��J�h)O�M�c�ct��ʍt��K��Z��}��J�?}��?��i'�%����4�` �GgkYL�@p:�Q�5{mF1��/���B�ڌ�4��P�cU�99AX|�,č��$4	-!\�<���A����xg}�-Ɵ���s�0ϸ��9�QK�\��G��/��r�O|"���)��;�C.ڿMyE�-�6f������o, ^���
c����7�;���۷�{X$��q�S�ۥ1<��g����K�j��q�SB4�D��݅�>B�?굸¶t��Ն��5���]�.._�|=���k��L��oA�����>�e&��BW�R�V��[e ��RǫZ��f��l��� ��&�	%ߞ��^ܜ+����(�s � ������+v�j�9�q�r��P^��"�"� �oD��F3*I�ĕ�Ӊa%㟥�%9қ���ppG E�ޔ�,�C>�Į����:�)|=�4�;����d�N�PO���xQf_jW�!bE`|��#AT���h�*�X���[�L��F���_Ó`l��U�_�V��I���1����F���'K�U�ʿ.E��j{����V(>�
r3`�2	�U�[Va4����s�����MT�&�/��V1�aU��~�^�A����,�H�E���A���	�4j���["F?Ƥ��b�r��S�@�@q��ZT���� c�d:���##qE9�X�KLX&�x��>!����N� �\x�!H	/Ự���3��,��\�������<�X���pw]�˓^b�n5��-�"����q޲�6�����S�v�C�yƞ�:#\�����`�r���+sSi�k�""��rj66����������;���ME1������#G�w�;�ri�54Y~��+�'�쏏��h���2؁�v�\���/_���H~�)����o�`��?��iQ��ݻ�y,ekJ���u?&��>U��P��,�ޯ'>�m���/�R{A�gN�B�חv`~zq~�+зN,���P�FL6=w3� -&�KN<�7n&s1us��4L;[$b%
�L�0v���"�c�m�[C(��ܜ.�k�X�����%�f-��#_�-m���_�����k��]���v�#b(�	gD����E������D�������.ЙO��N�o���W�M*&��Ɣ�#]�``i�ܕ@��n7�\�@X�@/8�$�@��g+�_�ɝq�(���BWi�k�B�E�l7�?ǪC,�?,slx�n`��NQ�f<9~8��i	\�� jB?��\'E}�����1��tC�'�ʏ��'�S�$L�����u��h�K�.�ʾ��|����Oic�_�zw3�9fp3?���"�W�n���ڌ�aM�F��_��^Am0�aTKػqr��.s�[�'�<Z���\�K*���I}��}�CZ����q�#�U���(J�#�+˯��������� [�!mAw��W�Q�Չk�\*ԀD-rt�nNRб}EC)�}Zd�D�!��6��#��\ԹYgQ���ռ�����5��j��=j�o%�1�*�:����j�n��.�r1�\�#�d���Yzj���Ӣڞ[� �"�D���	 B4v�6ʵES8ģ�Ua���W5X+�h@K��?����qr<o��꩔��$�ȤJQ�?��2�/#�h>	S\�:9�j��U�������;ù]�~����v~U���u�w`S� fH�L�źA|����,�?˕.'�S���h|w� j��^*Pn�G�Ʊq�h/'���\�$t"��k1���0`�ota���^s"A�{�u�0O��gS��,$�$�̿�(8���C=Չ�bYN�8�"���P$����w��ܸV�$[��x���Rq���ԝ�4�b���qDك�čr0�CJ}+dy�a��8�Pq����T���/�g(/G�!"�� 2�h�~va�bj������������QJ�^~I>�{/ �mpB�������Ïoy����}=�-�%)���P��S��Tq��~����1X:(�e��2PhZ^9J*���A�?.m���a��]�z�~�H?�#?�F�����{˵�)�����+�#N3�7�{�u�Y�?}<����������N'^y	���M7z�"�ƛpZ$�ݑR8l7������\k��=�7x�s�Xa�/�R/vrx�\\�c����<��C�A�7ݻ��ɧ����?���|�ҡo@P�	�������������i&�'?�l����]��{�+z��s��PZ\��VR�<�P.`�<
�&T��k�Yb�@cR	fk���g$Ehn:V��N���c�9@�e���n��oZ�
���9�x����.��4�%���9�_�,W���3��m�$�H�s=?�'�̽���׶h8)f����9���j�TѻgGoY����Y��e1����!������.����i�rT�~���?���((c���͝��㬝F�f��o2!vy �/6��!;�:�` �C���e���j��锛ʄ�K�L��Ķ��u�&�.��C���yP��h=�挥�h({��z�2sN ;��
~GϡU���ɮ �@P��b��:92�Bې�B���ǁ%�堍u���嫒�+$��Ǳ�K��w�Y��B#b�^u��E��z�g��;��57�l�FY��%���A%#�03%4���թ��wF�����Og���k�����x�\;������.�[<����u;�(��QH�Zݲ�d{Xު2fj�1�lZ=�S-B�������=b��ڨp�G��V.ջQsXN��?{��IKF8�"�O_���ek<P�yݡ�Ά���_rR�4���"V�"����������*|O7�<w�܉���QB���2Ak8<����6�؀���ֻ^�����L2�ᇍ��d@(���F�s�9�~���w����  @ IDATI�m�|��O�|��ԩ�S�t�J$�2IJY�)a�L����2V�=�<�i�i��"}������j�	7�ܫ��BZ�/'������g٪hK (@׿l���Q�L��@7�Y��JJ�"�T'V�m�zc
�΂aZ�q�u�:�w���1�͔�����~�L�W�5yӌx��Ӽ���[$��3(�>Xx.f�m-8�E��$��qLd@���l}P:a�P����믿I@C��%md��=4��_�'=����Zu�:�qB�P�8�������}m�����7G�s
i�d0av�垥?��Y���BU4���C��+2I���_m��{-��>��}i�3�u�����_�j�^��4�8���U�?��4s�H��/ds�����Կa(����1m���춷�;�s _{�����a�VΒ¨-�q��7��0�v����X����>�V�n]��ǔ°a�O��JG�M���ϧ�n��l�-0e���w}�H��l�@;Od�>����oHo��g�V?��OUn��7��4����TZ��+��r�*�+��x ��?�:vU�?a���K�����C���3v[v����z-�<�o_���r��C��k{�"s#\��2L���`�J<���g?�U����_��V�+;)���&p)�v�����x9X����[�O�Ps|��$�p�Α��_4���EP���!��,���5WV��^�J�*�}�}��b-�ex/���eXy��[~=;�$�3�*�utD��� `s�pc�i�(�ܤ�U�UD�u�"���+��lP?�P�x�J ����F)��Ml^&[Lc`�md8�޸�CBNc8�o�4�T�����6#�;㌺����+ �0���H\�Podn\�7����?��G.�Lt��+
����!���'C��v���;���+򩶯Hm���%f�-��Vm����Y��
���U���e��W)9j`֌�����hJ<ȷ"�H�V~dT�U}\��ʯY�*�ee��ʻ_�o>G������K��#�����t���ք���_����ߋ��^~5�[m���k�}>?�������3�{Z��O�Ze:�ĳ�*�ņî�I1���� Av��FF��)ĳF�1Q'���x��L�e�#o&��v�� �V��k����Ǉ�+`	;]��ܢ���L9���D�ݺX/˃���9���;yr!MNM����P]�>�qh�^r�֡���ۄa���̳[
��LTA���Dt�r2a^B��Ŕh5hk�l�%Y�Qⶤ����ٜ�^�N�	 .م�!p[=B�a�a���=p��7]ɖ�v�ׂDϭ��z%�����-K��������}�w��?�0��@��w5=�?�����Q��;��c�49:��L��S�J������%ʘc��EY��?�xIc3܂���W��������vuu���ۿM��{o�k��Fz���dz��G�vnN�m�����}�y{���]ٛ��?ӣ~/��
S�go}<5�G���=���2�x��6��Kf撹�I�O�<�c�n�} g�N�H-��3L3�|�'?�����X�w�������f;7mH��^���{Gz�Ͼ>=��}idb$�o�Jzۛ&��8�Ν�JC0��_���;���y���n����K1�2�H�$�J �|D��#�����<�V0��?i[�ձ <U��O{�R8���J����U�������d`�Lk8��_��_);�W��}l��� �ٓ�D �H<{��Sɦ�x�r���Y�2.�$��M�����F/va�7���ڰ��}/�2����<�x���[��{���_��/�Ώc^H?��E��+^�I�
)�\9R[�����le�����n�N��7M�+%��ч��#	�S�e?3������%=߂�tlUҤ�R���\AQ^�_���]+��m9s]Qd�baa�dKj��(���cGo-_���Rs�	�x�h�Z@#vVE0	�s�V�&�Zk	���`�2L,
�
�w�3���02 [�H�t��3��!U"+k��+�ek3��Pp�:J������e�s��G\^eX�w�⟍�ӹW����W����W�<�]Z�,���6�(�\z��tU-��v�E�}sv<Lg^^��!�r���^�Ii<UC��ki���j�^}#�i����[8�Z<��_�\�S�s(��nQ��/�7��e�?8�^�
�U��w����r �JtdH����3���c�}�lD'lX�~�2Y�rwA�!�1�Z�L�YɌ�Wؓ�ZxЖ���.N 2Bx��Y�&
!�"�o��e5\Y[�KF��a�0��l-�u�lA%��h��n6f�<��u�⒠=۾}'�V����*��ҋ�1Q0'��i����D���.~D�e���Lxl�O�����F��wmڒ}�CI��B�9�q;���ZO}���ó�2��I�f1�85������񑼩��S��#mYW��!��᳇a�I&8�b<�H-i �,��c�O�;v^�8��K�&n۶-�u�����`��a���y���9�ud���]H����lz��#u8������@zr�#���K��|��C�J��+�ٶ�/L?~0}�[_M�z�$�w�GP��tfr2bqN���d���L`5�D�ר��i/mj����Kq�2�Ծa8�޶=[n�dzd��;n�2��H����j��G?�.�ޓ�y������F���ӛ��[�o���c��D�쵷����wٵ9C��?����;x�[��Y��X_��Kݩ3�a�"��6��0���
�le&0�l��F�žZ�\W&���8��2L�w��P����H<�7�������F��[��AVt�S��`l�q��;�Bj����=�H�إG{�W��T��F.X%q"����6�T`cC��Ƴ^�w�ãM-��ӓ�q��R�q~���ҷ��e����ʫ������;���hŊM��Q�g�1�>�e)H�3-��'bHNM�%�Eap���qQ��BG>0���/�p��U�@$�ᑡ�ܪٛ]A�}��E�r�wv���c�V����!��Q�F X
Jt���[@��E�e#"U'�/�Gm�^�ՎX��خ�x@5��s'�W�p%d�����$��۬[Q͵j��eM���n�q'a���=���'��z7̫|/ފ�%t�}�����k���k�Uj���甿�0��.A*	9� S��]�U�?�l�2��o�������I_���2����&?'�a�������(���h2��)xv���B֋ _f����Z���P�e�'��1��r�	�+R�0]A�˴��f\֡$�� ���6�z`��v���<��և2C��ؼ�hR5;��y���5Ұ�'\Q�˘-�hյ��U_��}��6j/v��7��q9$�;�������
_�3V��y���/��~��`�N#S
��2���܈M�r�͑=v0{𑃩��'�E��8=��K�S{A�4����#/��L�)J�p�&��/�H"E@�`�6��([f�^D�O6��׏��|��F��k﵊�%ڰ1��7����?�mݺ�*��8�c]��P�G������+��򲗥/}���8�����![�i���O��U�Fa�&q71�1t��}��g���x{�0󅴣�3�S:�u_��Kn/�_����&�unZ�Q,S�M���t�G���}8e�?y,=��D�r���ء���^�K��ǟ��_�!��<2���\�,(2�"�PYv�:@F{��"��� �v,�{zD�a�6�?�ˠ��%T��#ߡ�p��Y����"���NV�n�O?����p��ic��╰g�/�c��� �i�I��Q�3��J�&v��w���y�`��"C�'���˵;�V�R�8�b{�_�=�mq��Z��c�
��V��7�\���nX�U�/��[m:�M�LW<�G<�̿����/�M_�}���|�� x"9}���ˁp�*�z즦V��cĚ��bڢ���ɐ�Ad.T���o�5l�y:X�԰�h%o�Q�蔲���Q���/�F��-:�:3�d�]O�T��b�b=�|E��f��M%]�1VڮrD�j�����%�U��VT�9�*��������F}C#�ɥ�����7��B�@�j 
V�5�U��<)%�û/JM�w�թ�6P�q�!���F�Y�S���(���Lw�p�wƵ���'��U����W_,�ٮ���W��De�jSb���#c�W���Gy�2�$ͤm�	Q�������(���i#}��'�D%�g����" �}�k1��qqQ�2�Z�����v���,��v-�y��1�2��pG�"�L_ԕ��Y}��_��3�n�rNt_]]d!�BB�"V����mz�?��"8sq���G���p���^�_�Q��8/�S�gɬD�2����F[�J��y�U��D/��DQ��>l�L��5r2RE���Ԟ}8����5�?NL3?�|��w+�G������hǙ3��C����ںٵ���]bP\�?��`+�R���E?	~�b
�����n`������ߗ^�/H���7��}�+���w]v�����OQ�T���uz��ߕ��@zŏ�DZE��܁a7V���M�GX$&=8��aȾ��2O����s��.,.F�0G0H@�pg�3�0��?m2�J��e��Ǚe[r��e���m߱���#��}g�����������l�f+;��grf�lWf�<p��4;	��eo`��,B��i�|Twa*L\m66�xj©�t����i�ӧ�9:dSz�y��Y䁽�S[��42S���_��F��;��6u�#���1�����+���\��`,5ʞ�����T��w\�Bv�M/���O-,�e��V�Ra�Q�/��
:�|��⁧Q�`�������-q�t3�����G�ꄱv�͸�� m]��	�P�GmO�/8��v�uE��18ze}�.u�҆i���c�U���7�|�sTu�3��QU��f������g��i^���c�ǒ9���746M㲉M�agCƎ�8w�k����7��T��w�}�[�lT�k�2~y��������_+���N0 ���{~�sp,5K����NNe��p��P=�}��7kd�����2
�Î ��ne�3��������I\2dB����#�U�Y	s�b?��Gh�f�r�"[� {R�O̽�T�"�ܘ�G���qG4� 
X��ګh��T���"s3!����GB#��8E�XEL��g�K ��lT7W��J��A���~�I
���:�����E������i�"�/��|hoı�E��,ƅ�?s����o�q���k���z�����w����0'?:�����x,�h*�h�I��T�����"����I��pr:�]�Z{Et?�i#�j��[y7�(��ըq{�|Ϗ�l�"���Ϲ�$���\����p`�N��ɚ�?�nDq�_uq��`N-K�pk.��L���&��?)ϴ0*!�G���yZ�O0S���oz�E~�=�a�I&��!���Ɨ���D}y�a�R�������7�9Sy�gH�[ۻ�-;wq�iK0]2�F:Cf��bg��k���<�.�0�J/�^p���I_���6�+w� y���!iP���2;�a�8�q\����.�,q�m�ڟ{uڼec���{�m�'��_��3ip}w���5;zt&]t���ӟ�t���|u6��Ѻ��iiF�a�N~zt��6$�i���2�l�瑖`|K���!�b�U:�n��^�����}Ѯ^��Y��8����'K�{��o|����ړn������-���?�\�e*�I�"���D1��;��]ѵ,�p�+3̰r�I�a��n;��KM�_���ŗ���"n�a���+��W~t�L�e`#�[[:��t|����;��[{��9v�-e����3�Ç�`c��$���C�}ct�x>�<��R�$����	��Tעg��Pk!=�v�_I?��h���+(�Y\<	76Xp�?
51} �$»pU	�l�x����@A���?�?�x5���G���P�S�q���%qGI�jw瓦Vjԯ.(�?�詓�^`�
c�8�v;��ul�jg��B<$n�8��o��w\��Ŏ苵g����{��gJoؿv��Y�l��˨��7����T��I����8	� dͭ8����,�p��30���H���WM���(��	`�1��NL�ɒ J����-c}�,�w�H�F@�qcx$����\����ON���2f{f�s2�5�g� ���Z�P�e�2[����`}���q+���#"	b`����I(*	1��S��͜�4b>���ՠ��<b�E8�32��a�̙��"�F��3X=_5y��|� I�N�0�|5# ��g������5�֎,�N �h_��dj+�碭��k�o�8�ǭ�S��� #9EIv2�#s'��յ"=��h���~�VL`��,�-�"�pެg���b 61�#���z[O ���-�8e�"UъjX1!�!ʯ��Z<�L�2��^�i�!^^�+��ᾗ�
X-c�2�=��Lh���3�4"�i���L�f��:|�"�I\e�,IR�!!�;N�7_�`$��``$�~Wbóy��My���H���P�Q�a���ʖUMgpن��
;&%K+L�Hd=C�6�F�L�J`r�-�c�'B��yTJFV�6���-�]�>�*	�--m�3x�2��	��0���\�p�k�B�����������|�g�K���Q}�囍Dt$�����曯M?�c�qtFb�?�_t�Ut5�[sÐ�ڶ��0�E��H3c#�P���s���{����!aa�(���ŶrD��嬩�u�t6����{�������8�"� �L��=��
#����P���n�Ẵa� Fޏa(����dG��w����u
�ڂ��`j!3=����k���Yf�q�?��G
�
S����� �6�~��� ���i�EBCg[>�0�5���麒�:6����NG��B�a�������>|T�#�y��<�)oZi�X���G������A� �H���%-�*�0��B��P�Pr�M���]�x�Z{-��g�`���݄p����S�/�	����N��L�1������RP�u��ۛ��v�^��Ϝ:�:V	�ɕF1��70�m��a(�9�eݱ�TY��;9)c�d;y,"���S���va�3:�w�M���^�9E�m����:�U�\~�C^���h�U��ټ���[�g�\������/�_�S��;�#4ʖ�dXUҤYViM0H"�:Zw-������yz=���]��+G���E "
�q'�89Mr�Z'u���)}/ɌyDÀ� �h��n�ͦ0,���0D�r$,���j�Hl! 0�e�QT���9��=.�t�
�.0���s��	`�����
.^
�P������͆��L��M��eqlq峧q�@?�q���(��?��X|8�s�Y����`ES��q��M��D�b�i���Է�6$�v���mB�2�ٮ�b\j"ET)#P�� 8Db�T$�1�h�I!�J�|�!<2�L�U�R�������+z��1�ع���緡�=�J	�ߣXK.���l�ʼ���̢���{��iq�1)��:�g��T5�-8����r��\A�e$`��5���J0%��e��eن�\��O�2�խ�*2�� ��O����|�S�K�eؔ�=V��_�W�7LO��}��G>��I��Uz�8@���*'vo�c+��Q��#&'��٩Ԇ��s��ky�h������0ơ�K��!a[�}��&ǘ)�������pѷ����mSC�f���m��M6�J���?����[��6T[��ڕ��n����hk2�m�~Qz��i�é��?ڿ4���
{��`�
�2��ܴ��.��� ]���*�F�
M0.M̢��wȜ���`�93,گ�ұ�[�;�<G�M��{dD��y�l����ӠU��	�4�N'�`�J#���wg^#��`<Y�(��	Ծ�*��t �5��j�I���R��`�EE\�b��L씎Φ#{�B����Fl��aB��{�+�Aj�t��e|BFF�fSs��
��UvS����]j��0��H���,�57�Nt	5R�@�#H�I"UsI��Ԣ|
864p��O�8v��i��o��T�>�0�5
|	���$L�w��{m����kɶnޒ��◄y�*���1T�»$_��&�xu�&���}6=�Q6���콘۰3C{�Q���$���J^wH���9\v���*:1攧}+��ڴ�K�;q"����OmX��l��^{զ�-�'�ǢLYK�i�@�x� �vK�ȴ
bM�:�Ϗ�ʶ����ɲ����ٞ�̏�4c ,pT0<8�^N�H=ae�e+Ksk�T�X��^TN������ K,`�A��K���ӺΖ(~AJ�:�WQ�U�|�ڵSs�+��Z2iy�Sd�@ T!���0��C"f��#�o��gB��i���
��/+L
�1�{���0��ca�Ԟ �Bۦ
}���G��
iB"-i�����z#T��X�r�ȅB������! �'���ABy�:�n�-���[M\"T	E�GM^��;6�'kBH-�{b !���D�3�M �h`%ן<�]�r����e��:;H�{Y�(�@j�
F5�q��N�URMD#X�\���P��������~N`��LS�˸���O[Ə6[]�aq3��&���K�,au�������A��B",���?��ܫJԣ,�s�n6'JW�8�3o�\��_����֟��+
%�	���c��[��ƨ���U����0(&o|�u�|�B��8;vl�	>���j '}0iW��@Q�|Ϟ=Y��[�&Zq�;|ό�S����5�����Zf+���������]]����C3ᔋ0�	�I�GspHR�����$R�Ʀ���Dv�?;��Chvt25��XDR���G���&t�+��݌�nW���I'�m��BM�@�V�����:��e��u��[�����G$� ���y���'��͛��Yv��Q c�����aϥ�㕩��u���_ど,p��=��1��y�UQ6�NlgFH�����N���)D���Z4�.�J��4N�A~�tQ"�ڔz֯c�o���G��{u��&���+���hfk�=�!�jf�.+*q�ŸS��4v�շ�S�H�1T�j�g���c�$=�V	{H��^���%�� �PdA��Ob���y.d�C-L��.\� .��.F<.�ԾG�!S�(�Sv�N�/e]��%,��5������w(��{��;�Ǝ>����RL��Ƒ.������lnv!�gG�E�]٣�0���oe[��Rc�����t�J�\=. ��
3݋����/ ��@]�D����x��Α�.�u�N#��3^���B�W��4峟�<�{m���i�8�)ý��U~=[���3���iYsein�XZ���/R=�χ�Z�����lg��	v8i�z-7.{��g@W�����c�ދh�$&P�<xNZ3,�Z��",z״�p�y�.�N�3p�D���qj��� 3��
����)��0�����F!T�����_�T͍�)�)"{�gz���V!b��pm!!ApF�E	���X\��T0QK����]�k�U�.(e䧇W��Y-��6�^�C'�6Oe�4�;��7YV�I����AT��ui&ѫ��׼�-��]g��RD��E,����T�(����.'�UA��D'�̍
J;e0�~��
Da�Ps�/XV�r�\a����ß��%���s�����mlNp����[�k^�϶���ܯ��+��<�ު�ֆ�X���4�Zl)¾pہ�2G�+Ҋ8Fǣ( ����P�D����L6W�Cgjj�m���260=~_�)�H�UO��P&JS�&�`Ԝ��H.�K�o�ͫ�Ck+No��qE��,�,-��&�?veɰ-V�ALՇ��۷e�4�a��U�q&�>\Uk�!���d�Ū��X�e�h��%��B�f[����L����O�l�Q��̓��Qw|��ϲ�?�9m�����3%Kq��yP��+R�Ԁ�9�^FU41=��d�����&'O�Y��$�Nf�\wq=ώ���
����(�7��`�2����c�Ԥ�ML'�q0���؅^Ff2�R	��RG��?���:�ԍ7ވ��EH�p.�*���*}���@0%,X[;;V�*c�'�*�ܴ�d.�Ǟ��r��}���=V�d.A�08�`h���!iK�������4��i�Vi*lk�(�x�~.���.㕻�'���uj�� H�X���1���V62@Ga���E)�U;����C-��*�}�ܮ�8ˉA�S|���)���U`Yݜ]�#��Ip��x)P�0S�+�y�0�1pE)��ή�8�m˖-|g�#���S0����$	�`ͱiCi!VQ�J�1A<��Kӎ��9p�$F���nǱ��S=�&�nH�6c~�[v�8t��)p���1T}����3+��e�W"�+�B$�C�+4��?���_r�_|�eC�w�g���N����^��g�r�e5�t����g�d�a���Eia�,\�N&�
;r,��#=�X�ӿ�t>�R;@�O�zR����d�x��<;����� ^ ��仕�g�˻��Xf�㯏�$׀�t�s��ͬ����3`�L,�vJ��O�"#�ɹW�4��X)X���2��̠�Gҁ�Y��'~��c��(*��PY ���81�U�@�OXt���;vTU ƍr,18 ����)���euƪ�����d�DD^:��R�f`R
�P�#aJȁ����"�Te��V��y��������E���W�g�!�\�P	��QJ���*��!�2�1t�te�;ZVuKzd�p4��f@q��T�,UE1r�s�|XW���K�\�>��KԒ������R=�h��7ғe�F z�U�qT������:����2�a��e�k�i'/k�~+�Ĥ�{�}!1]� 룧��Ɏ^Qj###3�Ѳc.��;�P;��%�������s���|̘'�02E��]�0�W�l�G���V�C�.��-�*3�c��ݲk��Q�͆�m�u��YI��Q�e�����L��D�ri�*u <�U��y:z#߭}���Zٖ���񃧐 5�W<�9Y+���G�4&�^�:��!��+���y�[�49	\�/�l�b���|��Ks�d��_촠G I��o|3}�_jnS�ʶ����X����yÓ$j Tt��r, :jc=}�C_[1,�K#�W\v�%��W\����*S2�-���ɱ�C=���@ںm3�rܝv\��
r8,��@�~�O?�mg��f����݉���i¡C����� �RڲuK��>ҋ[^��i��z����z�zY�!��!f�]e��T�d!x�Ҁ�������Aa�0�oI�v��
��qcjf�\���s��#-kJ��O��IM�CҩIav�e�>�u�j[[+����4Gn��2uåQ�*4���C�Q�F�qvlKI��e�C,�ɭH2Q���&p-$�)=�đ$��~��'4x"( ��Wl$.�2�>��PO�ʼV�I�i2��Xܥ��Gj'������[�暫*��jOO�:�Y�_b~_圶=
��I�������u�+��#汰s�l���Q��)v�-��mbW��v6��(*�饺�i�a\?.� � �qYo;����l���Խ��.X�Wgg�q�S�?A�X̓|
ҿ�]ݡ��'����B��
��bu�2�547�O+wL.�B���%���c������Ќz�H=����xbj�:ʯF/h�,<8���ZOEc�$^.�S!H��{:���6Nn������Ճ�H��.m�:*3�`�H�pqI���W&/�*��8!٤`8V�8V4����[��q#��.|�sg� ��%�2�Z�5i�����ceP i�b�y
˪�k�q���]~��@0��W׳�����8�nh5S�ؤv�!w[,���/�>h5�|vl��4�d�x�a��0�jl���Y�u�`ѭ�9S:"��9�P}?�`�0��} �~S3�@E��[�
��/V�n���fhs{V��₠�\��^żhY�}\��ՠ�o1�V���s��] TT*��|*���?;U �97�lL�*��[�k�N&�?A��*٠�10�E�4͢�-��l
+���.�Z֭�^X���ϵ����6�>����紿�Xs��Z~�G�#�����Ԣ�G!�X; �@b+V`��@Jʸ�XG���̳��+A�m.�(�(ƂxLHJ�b ϊj2�q6��̑�HY���F�J��NQ%><�@oWƨ�nF�Mܨ�:�c�T18!��扬�B��?��8���P���铡�#�ph)%���H�U���B;�wH��"r!�!t�GS`Ů��y�+�S�l��@,X�)���L1�^�@�(p���~$G�5�V�b��{0�� X��%ҏ��s��XT5�7�8(���}T+L�O��ǳG{0=��#����vn����~,���Зi۶m�?�����}'[ЧP���C��$-#Fݲ��O����ǎQG�xw<�@����Jz��r��鳟�l�����׽ [׻>=���U�q�Zck[�xzbϓi�ާR�������8'i"XpܧqL��了`��(蕾��?�ദ�����<42:�wv�g]�m�8~"=|4���&�T��g-���Ң�<ajLo;~--��KS��Piț�9y�V#ަ�U�$�����BT�l��E�,�	���	A{f7I/�7	Tql�XTeEC-C"<�G�e��s&��ѐ�/���Y��0�7�(v�)����M�[�V�w��C��oCx�t�ȑ4;��s�;8>ϑc�Qf�JQ����G�?a�ς 	�k�ļ��!FTM���Im�������N�4�5�[�/$���}����.މSІ�}���������u��1�A�Fw���g%p���bi`~���0���a:B �R��H�+��wJ'��Ho�Ӣ},,�`㈘�%$��0CJ����Kp1�}�8��uX�_A��z�ӊ�3^1x�sH;��Q]Gt�g�'�v:����v'����3���O�҆�l�� 8Į�����r�x/��I�2p���E�9�a��s��#�̕���Z�L��2�[i���J#���Yq!��>���uq�={ߢW٥�����G�6Q���X��a9�xͶt���F�lZ�J�zV=XY�c�HΡ�;�,=�*��=����J�Fv^� 4�l���魿�v�O1"�I�8���7�6���x�g%�M��r}~��H����L��]�g��M��O���ȭ��??��{�Q�f�U���J�`>}��܎(_�I%R����4 ���?ެ�%;�(����N��W���F�X�w���v�l
��@��F&4H��]�9� z0��Y3���c_��++�l46��~��Xj�.`��Y{e!��+8mAu�ű�K�lXH�GN���N��9���nE��!�^F5���<1Y�N=���ҵ;���W\�z�w�V�C-޳9��50�#�pb=
��Y�@�L�,I�M�^�R �D&�p/�Rpf��+`��Y<,69�������+bk2F��&�2���w5;�PŘl�@�(�������3����H"Ԓ@�b}Tt�Dy5H]K3���&Q�snu�p�-�3ϸ5��QZ����%���xIW!B<�W)QCH�$�2���+���UN0W����>��Fad��>|xH��fH7����Yn��N�Z�W�a̚`�܉�|HVPo���8�s�Z`8�(DC�6b�����d�n�^�Q�@?��#����4�-�f��:bP[mH٢�3�gɄ
	u�jۏh?�6c����m8�1A��R=��18H�^�%&��
��*a��96e|��i�C4�)�C\��
|�O����d���PY=sf?��c�w��4<Ԏ��-}���^��������O=ű������Z��!Aj�0�N$%�7so�yǎ���֭���s1�;�[�r0p辘��7��J���/����.���[���jK>Qٻg2��ȁ�ѿ�fv�%���,*���S�w^���6�ǉE�"v�J�/���p��{i�� !S`�9#�E��'޳��;��Qe��H���ebF��9O�^�ݍH啚�1�<��U1��1C���0>m�~� �e� )Kt/A�� �H����1��4�T��]�^� �(�7Hen����+N������K�d�A��i�	��H=�+ֿ��>��;�!�1Z��7�E&�[����y%�2��֧^�c!���@#qg�E��xH�`� �ԍ���;�1�^�F�ؿ~C6�B����s(3��f3�R8��X5���	�Y^=5���XZ!C�)�J��Aq�������ԅo��[��7O}뒛(L��)/�p�J������p�w$� j�WW�����E����l�F�6��?x��Y�e���d���}l|�����H����@��� &*��`�
�F��$DH��Ū͆O��p5>:���uiV���;��I���L��Y2�d�(��d�蔘��C}_���-����x�A(�2T/+l6ލ�UY^�]=am4P]x��9D���C�.D%�Pk]"�P�Ydu�p�a��S��],bP�����?�?us�ݏ��Nw�m�p�V?[�9
�*�fW��1&#%s���K�ɍ[�M�^���o�.צ���[�%7�G+�!�1�Y���4�!�u�/�|�Ut��i����#���(���ҍ��ͩ[�y{�6$v���~�_������u�]�n}�-9�R�{�ե�|�#�w�sR{#^zANfKΈBV�D����n+�Ӻ�y��`�@T���3��HP�QE��N�0J} �����uW]����_�n�~��66�@A D�孎Q�?����w>t0;2v:��mϧ� ]M�L֍0J�?���/Io�O?���Re�������{8�i�ܛ`��Dv#1�R%���Q9�p�����?e����_�y �ٽ�g-��Z�Ώw�{D`.��_-�k�G9	eqQ��/�z�_��{�	�kH��3���U����C�Q[�!�A�$��*5��8yI?̫Xɵ���%q�!�%2g��ɔ�q��e;�ȜI�ʺ����`��,YG�%6��C�g]5��x��lg�9u�D�w��lu�xG�i}��<ꦆ�V��/vZyDPh4���D��G�"P~T�h��
����E��s�2M2��8�P�g>���}�`�d�LyȊ���[�a��f��}{�7��MHeR���>�#���+�SLB���(���d�p]Α,Y/x�߄ѷ��'�x2$E����U���VN?��O�����즛nN�02��4.Q����w]�G�t�}a՛N�L�h����-�L���x�fR�p2�u�D38��	�Z3�&�{M-����<�)ƿ�#c�437�}�N��y8��d�...�	���.f��8�q�K<�ǘ��:� ����uK�Z1n��C���V�
,��B�waU�����+a���n�q�Ԑt���]D��dv�^�tA�d�3���0o��C�3� �Ќ�vv�~�ήj4	#��f��s���OrQ�G��Ql���Ǒ ��͆7mBu4��y���l0��9u������̍�m�lȐ۾�����U	�;v�tR��g�SI���1���b�tY�W�M�P���Ig`n*���1Z�8W0��E?J`r�Y���Ku��j8�b�����`�,��
5�e�]��13�����S^��H�����>�H]n�9�=�����/̚{zY�
�
�(52��;�P�
Y��.�GS��=U�  @ IDAT/�Q�Zh؄�����u0��+�5���(u̱�n�b���z�l4>�z��E��v.W	�����_qA���7�i~sgF�w��_����K����Ȼ��rY�#pI�_x0}���F @���O�}<��`�6�VR��w_�������b�K��= ���{oM���Up�)�QKW:߾����ǟ`�\IW^~E���6��.�Rv�.� �X��x��;���y<۱qC�����BAf�ν��5�y�ci�1l>د��Ґ�:{���t�sv���,���M�rc���tj�E�k�?��*k��8� $L���iFO1C8^���ÒX_����j��hL.��4"<������o�_��Wfoyí9��>p�}f�	���+��p��ozU��O����?I���6r� jn�=d���L��˯N����i��-�+l�O�l�Α����	$UZVhձ������ ��6^�\~+�X����ߟ�y���V�]��eԆCB��[ĵp�xL|��%�nmb�PQ�_m��w�2�G�Q2'�;��.OA��H[48��6F��2	J��8*A�� B{'a��(A��JZ@�m����&�0��3�0�@����+N����G�x�h�O�菹$ʚǮH�Ci6o�*��%�=}[�8�s��)$��D���&��|�!Tl�[�����J�0\�W��T��u��DDs��`����"ϡM��=�Fy$��I$>���q 2@��:abv�buz�j_�������v�H�~������ϧ�|���VK�V�~K���Q%��f�p�����>B�Ǣ�\::�ZTz��"X����SL*����]����#mKb��7���J��ؼn��i���ߑ�p�Tߪ�NB�n����4]	!�q'"�O�n@�Gr4��&�d�� ��U�%BC�g��Iv���#��,�]�TL��k�h��OT�`m������s�`��1���w���_R*A�	�x��̣DJct���B�z����ɀĐ��JA[pjI[�^�4����C�=�_���[�C��n >��ۚ����#�#�����L`�۰����!��D��XJ�6�K���9��2ܷ2�mt*��5ׇ��9>�������W{0o[��È������em)�N5��,�y�#W�%�"�ؽ{w��L�~�d�6mި=ۼys�qVZc�����&������q�0���;��m�������ו�x>0��n�b�v�ß�[~��"Q�܃�);蔴
.c!��~��F�x} ���s]b٩{�l88��Ѡ�n)mں%����N�BJ-��A�3�T	���Ab�$|Bm�/�M�
 .�5Bb�O���Dgm�@g��X�%�6c �� Dq]��ۥ$a�&�"r�a��/�D�����H��%BX��Յtr�T����ҁG������#�$�* ����#����T�;���W�~D�+����8zܼ�R�������^F�i��k��\������5���O_�?{���tǗ���Tɦق����K7��E���.�n�����@2�����ٛ��O��C�h��w��/�L�8s<����?~x4�h�Ŭ)�8��������7U^x�&�p�i;\��k?��y�og3#�SS��K:���O�D�E���2Y9&O�_wɡ7c2R��LեcbX�u�/��n��2M�&�S�]�W��=���̤��=������{YQ/��^ڕ���k�G?yGj[����ސ����^��M��%2gYE�>f�nГl]�v�.��v��]б����������j��>��"X��D�5qk�k��R���囿	�x�H%���O�g��C�G�<��N1_�`������� 8�G�H��Hk�x��U��C%�N� ��l|�A��J���Y�m���c�0?�!^L��X[g�~�
�q}����a�A�:w���DJ����Y`hxK��[W!������m��KnS���+!�Lh�?���n$�3�RƠ�WUZ�"M!h�5]�4(b�9��q��L��cO�&	0���a���8�����/���k�J5`F ��JȇE�K9�hY,�S+�3�'�H�?���铇b�y�[~��3����̇7l���:8�d4x����r�'��������p�8�7K���Ϝ>��� $t7^�b�z&�}y��˲7mM�~�~��&�.��+��W�z���m:�n#GZ��L� ����-i��9a�l��S�8�d�#v����%�v/!�&K�Y���s�T�ޭ^���W�M�}!�CY�	oE�5'm�<���"_�<$,��@�@��F>2;Q�_�Gc\���9VF�K�E�4�s�B��g�	ҡ�d�!�L�̄җ|b�T�����9�pGм#G��u�}����E�Y���??��w�c�S�ӕz�JH���C��^����¢���o�7m݈'�ٴ���{���3�l�hO{�:�f&6d�Hl�C���b�yA�Re��)N�o��F⭲3R��`PN; ��Ͽ�T-��!m������R!��z�n���ǣ],_z>��n��c;V�EڤT��*���4mx-�����j^�Q��m�P�?Ċ�'3�R0׭d��f�8`��"]c��������7=>����BD@�Ln\�B;L�����+ )� ���%|$n\պM��
[i��ɛ,�kyrc[(z��
�E�$jB[�U��-)����"��%�PeNg8ݼÍ
��������߸/��%H^���x�w��Ҷ���F��E���6\�Wں!ty�8q8䡇�[o��b*�/�"��&{������/ߓz�_�����FUo�˧g��?��?�M���������+Щ)���`���ҝ��������Hw>�$H�9�q��=?1���:���K���'�.�ޖ��8P��_���?����^���i�����+v�/޷=�0 �ɉ���j�~�L��*����9b:Ee7K�T�х���m8��Hz�����Q��o����9ݳ�D޵n8����ǏI�|�K��?Lzt���m�����=���<�.ݵ+��7~)�v��zʁ�T7�4����^fg�V+ln��-.;�8e�����U�U_�n%L�~_{��f��յ���Z|�a���7�i�ڬ�W��]���W�;P�#�s��F3n���/+ǜe2�$��%8��ݱ�a(jƃ���ʍ�+�p���sa�-��A��K(�U��*�R�]���
>�ʯC4�F�`���J	��qG���Xς($Vf*�n��/��˧�'��9W��T.ڱ�e�g���a������_w�.MYoL~q,�R��q��(y �XX9�GV��:J[����u-��c����� �*DdӘ\4�1v��jfr*0b��q^����zζm �K�ҟ����[�9�m:����r�Y?�(Ϥ����>��lu�7�� �_��ײ]^�ϡ��~�N̗��,�d?9a��4�16v3*:�1�P�e<el��B(	�Q}wwwb���${�� �}��Cj�#v����km;kW�
6�
������̱q�6$���eF�Z'P��f�v�̳��ŷ���̒c�k�����Y�o��*n~-c��ށ�b�n����e�(R��!�����O��X�X�"� �W�g�c�i$;�YD^����3��)L�F��C�*:��b}�^�H=0�q;@������	>������B��H�n�w�L�7slKkG.n^q�s\�T����
���si��C�IT�`�p����.T*�]:@C����.WQyΆ4��Kv������Ԥ�pZ�ҊL�m �Z`<ꑎ�Ӱmfp�o�/}�K�����w�9{�u׵us����l㉓'�������D�W��s$�q���2�K7ȫ��șŹٹ��6�3����p������V�Й&`H{�ʁ��K0rT�^��.�G�k�d��e+�D�HO�=�% ���x��9%% <�$�;�@3p���@����N���b����#vByʅ���U����`(�`  �]�o�r3��K���G� ��*P��UV�(�+ � ީu��EV���(�ᰕ����E�\�4eGR���Ɂj�?�H���~Q����EN�,v�Ԧ��4?1�7b�7�^EG� �w^rY��^ėlE�D�ё)�G��U������Y��&rT$�zdh$�h"}�k��z��7TN.7�GG9���7M�p�0���w�Kox˻������K��!�b|`��㬠��aΨb���������t��$Mpi�.�'�+�����p�[�����Ȯ���b�����J����e�spe�AwЭvWt"c�l�J�$
����z����8K:�O�R߁�9������d����tϣ�����g3�q��axݺ�'��_y��M��7��s�B��^p�%��ߞnx���=XI#��EJ���$��AІ�GK�l,���0�#U1�)��U�l����e��{�p����e����4e��i����Y˯�iڸ���\���k�4!�
�eP4��	�$��:^1���Oܠ�0������A�l^���"�������z$6$Wi���ᦁP�3wˀ��m�	Md!�eپ��+*!�e��oN�U��0Z	(b��W.D�x�Ƿ���k���e�l��.�1g�'�T$9J��<�4'̋����<���:VL�"�¢���&������m��I3�9��U��j���fPk����&I��r�|��+X]��Rڻ����k_�J~���|��ާ�@�2�Ql��׼&��?� X�|:�AՓ�h�ȅ�/��%�6(V��Ӆw衡	��6�yK:�ǁu}�a�?�p�|qt�Cې,�[e~f#����QS����y6��"��4�EI����1R��v�	�� 7����l�J
����Ɍ� ���~3M��f^1 ���g�x�Jp���ȢR[-����;ֆ�Z\�i�l�I�g��.f%'��rK��'>&������	��u� �� p֩c�
�.�;�/prW�PHpg�9~fg����/}�+H�
���K�)��5UQx2_J�]����+���+gfg�MhM>��/�C�K�!�� !����Kw_�O��g���ζ���T�b$�,�:M�{n��B�ԍ��D���`�&j������5�\3��qhh�n-:��u���Žp`�)Ts�����ZZ[��AZ��$��ϛp*:���:>3�п87Պ�KP|��3	�'gf�a,�X tq�o��:�u�6v�-wt�O�a~a�[���8{ փ�O�>Հhy��C��i���.�(�:�c���[aA���;^�.�q��H��Q1g� N{gc�~xC��l��TA�`y�H	�e;� [�¢�9��l�. �*)�YP��:\���V�/@�wɅ߭.�Yc�;�0&C�����$!�&��2��&S�`�b��AM��\R��d��yP�v�Ͳ�uQ׀��:!Y��LI:Ɩ�&DƝ0{8:��7\���k~8{�[ߝ�<~*kl�CG���@�ق��R{F#m��/��?������R�t����J��iאF��[vd{N>��y��.氕����h�P�>�vtg�K"ٶ�����M�����N]ΦQF�n�8���Wҷ��X����!U&f�C�|%�"/���.���U���0Rv�����>��=i�)a��֍ V�Lw�	�U�g�6f�%��y�!���~._�\�J[/[��z��Js�p�փOf��SB��Xl�<���D��z"mXߝ����o�)]�}��F����C>��֜\Be*��`Bk+��h����n�^~γ��z���|"�+�eBQV�/�����}�s�exm>eX�"Z鳚(�1�Dy�Q�.]F�G;��&>"�,߸\f�� W�����o�q��K�t�@�C|��a��e���4�2+�w�r�|ËzŤ�j�	u�'�j�H飍����$j�v���~*?~�x�SI�$�����2�k����d֎��:�</�6@AB��C�G���<:�gB���X-:$Z�=\������UYR��(mqғ�;xp����=_MɎ�C<r���u{���kL�5��`�4�ް2������'a6�3�J#�W�����FuAA\��if���pe;Yk�ǎ`PO^��eƔ����8E���J�VӃӸO`b�>�M'GF����cA��K.��c]b�7�D��X,�f�B���E�+�P�#AY���j�v`���RўE�A:s��q|�M��0G�?]ΰ���πU��2h���AR���cl� ��+f)��@R������x�_Q��q��|�:V�AXd&-[��#���c�O%�PpBƻv����%�;�p�(p��=L?m���&�#�b)��Q�m��ż��	�4�ȴ�p6���O�Q��$��<��g؅m�������x��+_G���ξ��y<�?S�L]�7�Bv.kS"Ƒ>�{�O����_}�飧�����m��/���|���Q�_��c����<j����ڲ�g����i��G��X�nx��-�(�R~4	�h�����4���$@�=�(�G�y/p�G1�|1��10���s9��V]�7_9��!"n�PH&�HI�I�I��8C��W��~�(�Ѯ��!�)_"[��k��� b�"T�E�(�� dU=��
�>�U����Eo�Ei�Dט��
��� \�2Ҏ����gz
o���4�P�A+�ش�5��`F^�I���ٕ[Rz�-7g����C��/#魯�.�֒�������+nI7�x}x���_��������|!�ݏ]O��!��� Ω�Im=�?��t��6D����3x����z<�������0�M��
nEsA�;+�4:q5�D�<z�<Z�U�]�b~��ޝ���~�B9�	��s%���V�.Ꮯ�l�0D������sg�]a%�����Dv�-�E
�j5�����ew_zc:zj<�5"�0N��-�������;���Wf�N7��9�%�/�E�����To)u�/��.ߝv�X��=�>�v���#��y�OU}����y4�־�^������EB���� �j�5�},��w�j���ٮ�x��?�����"�j�`r�P�����9��5�/����x1��M�7e���D��,�x�)��I[��%�*�KL�cc	M�L99R��_(�Iл�����OIP��h���2�q���Vn���9�����4R �u��K�3�s��
�PUn��m۶�&I�2��ԾC��v�����3t;�g�����+�� CUCި�r�CJ�45��QG�+��%���)��=X�ńiVϱDe cp,i0��	�@�Y/ƨ�S�m�M��	�@�&�1��XĲͺr*_7�;��F���#e� �4�ۧ�s�Y�B�g_.��4�KSK�rb�#(�������vݪ�t,0��+�'vò˭9���9�b�pKrr�Iwv*�p呷b��T����!��T5�e�%谎1م\���c0�~(8p Ԣ����i�H��/@s�k������64Zg��h	�ǹ�HD�r�FF0�a����ʼ
~��x����k
#Y�"�]��s%*�^u�)�Q7,j�+�2Z��4�f@������O_��b�V��qaX�4�ARjx���wz���V!���1c�d�W�+c7��pHt7o�S=���]�	z8o���j�S_�j�v����-fM�G�H4`�e�Ѯ��GՑ���S����]}[�1<��ߨ��*�˻a\܊��^�O��-�k�:?���e~��/꣸X��q�\>�Q�{�q��{YwfNEy�Q@� ����s"��\���J�BA6�'�����p�6N+��zV� �q;n\|&�U ���1�݄��.ED� s
�"�}��Bb����()��P��	��q�1:u�B�$�4��Q�&p�H��U gzI(GtX;�W"ABv����q�P�u�u�K'Ʌ4�&?�����ǰ���MM(�R{�a�;��P5�ܐ~���gzɵWe��g�4�͟{��y��>4oo~틳\�+����?3���G�����5M>������{����}���E/����nO�w �a\�n� �O��+D�90]R�H��<8i�q���#��7\�.�@Gh��<hq�d�s˺|s��d�p52�8mle�[�y�Tj�2�q�*�8�����Ȫ���-upL��C� ~��|��*��P�e�a�J��-s�/�A{�LeY����>����/�R����W�;>��r���ly�t>ݢELH<�����vH���D���ǠGD"�?��4<{	���s.�6~���G�E~����e���՗2���2n�=0�(.���ʧI�z���&�X��U�h� H�%��x�'��G
X��5j)��؉���jK�%���'W%�2+V�ի���4�0�$��K�T�<���Ŕn�3��
����b�q���8�$a'����κ�`9�`V�-�Ζ�2��U�i�ɱ;���.��aԳ`��/���<�]~��vf##x�m�Ά|;�<1���t�*�O0��)�6����y՞jE���\/����:
@eׯqH�^W��lQ���1����3���4�����G��4��e�ˊ`��1s��<n��wF��w|�{����ե��bG�C���.\��u@lD�
�7��M�D��:k�Yv^1"0f�3�w%$�'��H��?&�	�S@l�h��Yi�6OpH��Q�LO,���Qe��a4A����lh`�蕍�8�/j�J<eD�PU�&fS��#���"���D�M6���s�N��LH>�s��#�hc��@%���'#��kZ "?�����J�'z6�1&Y�7�E���YB&�q�qj� ��Ӕ�I~9ޘ�ر��rA�R�p��1wq����"c�a*Tڝ0�H�s0Kl����.��v���I����'hә�C�lߙ�<�/�7Q�+�w���ӳ�XfY��`ފ��M;�{�0�[	�*D��
Rɾ����NM-��U���b����.*�򹼗��2Mm�g{6ݳ}3�̫̿�[����{��6������O��DۀD�]Ļ�$(�ΐ�b�  (O�.�`G�]/L���n�Ȃl�<1������ŀ)B!W��0PG* )�������`A]�4��f�
F?�ڋ8xS�u&������3��� �E�\�rP��!�A����-c�;� I���fU�� )A�9�DM��MgY���8I�����Ƿ:ҋ��;���g�z���׺=mܚ����?�p�������;��k����k�O��PMQ�^>�]y��Cq�#S�?����{�ϻ��r�7�HW^�������7�yڼ��� ީC���b5�a%'�������<֥$[��eG����|u�h6v��������q���Rv�=w�s����v=�ߛp��(&�������,+��y+窮�i:L��f���a@q�%�?E"WY��"��S��U�5�	YI&%38y�'O����ꮮ��{���{��)f0|��n�[��s�=���<�9OD�if�~�^���Ew����^i��`w�JZ�S���:w!_vp+�����\b���Gtڂ�_O�Ƭ�T�(�/�5S�$�m@�n�6P������Bu	r
�N�_%Vr9�W�4�K1��c|�6��ּ�=]�����]����oTe����<�ӗ�#�a��F(t?.,��@���J4� ��Iߏ�G��缇�0��4<s��Jy����aq�?p�:�Tq�(7����:�U�Յ�2�t���PK�c�ĉ�4L������bc@2[�BdHL�6�/�! ���_j��x8�E.����N��B�<�mݥ���f؀�I�e 8�$4�1DO�E���И��
Xvq��5��m�%��<	ދ�V��a����L��575t':$�@�}"?�rr���v7�$���9R��Q��K.ٟ��oB���t�?}9}�?������8.ܶNf���q,U�F���p�=��(8�z�7��+8N�f�u�Y�i�]q��p����<t�`:�ؑ\\��^����FEw�>�PB�
Q,\/�Gѿ{o�@��pq9oݱU�Gz㡨��T�Ze���:�����e�M1g����.l�Wn�c��A��x�+�]��Xa�Y���,N��X��C��	��r��ʿN�����ŚD�q��� �(vB��'��ʌ���]vY��k�K*CK�3os7�%����I5�t��7ɴ`�u:��9"����x�mQ��Y( 2��ڝ=��[��856����g����(��q^wW����S�$�����ÄI�������T}A3lnU�y�|]>�������[���<�;UzUZ�������������^���?jڗS���R�0,0���!�UA(ɶU�!!unt���À���0%�F=v����R�p&��<�.\mv+f�9�J
���I�JSL:�5�!Z�t��޷�u�%H �!ic!���w�HI(�|w 4FL�`�E�<T���D�:�=�5�n�tv:�Ҫ�>X)�1/ބb����Z�n�n��xJ���-���O�}ٜ.{�v���Wݘ~�]��VϤ���o��3�Cx5�L��ܫ���^���o峿��O�����.\��?|y:���"�M����	E�F�$�>������}_L=Dtn#J6����X-ܾ9��O~�x1. 0��ut���m�v��ظ���0G��5���=�d9;?��.ƣ=&�v��Ʉb8�+ ��4	;~x��X�͝xy����Ա���q����GSkO-l�*&	�Z�Π�'����+��EZ��`��C,�Ĥ��� Ԋ%���j�V�R%tE*`��H�1#�����h<X߅���yu���սy7�Ϟ.��<�ќ�|�\����O�6M8v��/�@���,�"X�s�L��Bn�D��@T�t��pZ����{���`wĎ��Mq����ubG�Q3<�aV+���Yc&��;L1�i�Qs��
�vg�%<��c�2��<M}o���P>�=s.6z.��p�����7���Ŋ`]���#�U�pb�bt5�!���,(����E��bk��ie�g{�Sv>�ܩn"�
,�G�Ƃp���N��K��`��``<џ?���h�'��yc�f�����6%(]�9\���;@���2�0�~�'�sz�{�b�x�n]����CL������s���Ɏ.�(cɁ5(8pD/��3��`�/�%�ݍ�/mڵkG>����\��Oi������33i��va��Z�c���p*��GZ��,ǯ�(m�
	n��:H~{�M��	�Y���UXC�������V��1[����:�k�CⴈkN��O�#&�V�#�!F�=��� �E���5�;�@�G�.}�M땵��6���j�ݔ�y��E����b	�0'�$}z�1���2�*���bɩ�K��W;�u�ܸ�>�2L�>�$xU�߱{O~]/u<5ݟa�193�o��y�b��]�?����c�(���0�xRo�(1��wC���G�N[{:;��n�lϮ���i3�mt�k�g��|_���|�n����xo~Ӫ���W�O��z��_�{�us��u���7o�*�*���n��C0��B"���z�����X�9T9���t���u���.��1�ESO�X# �L�4�܌~"V�C��xF�R�����l��*X3	y� ��=a���"B�Jv/��A-mZ��~���l�ܜ�JK�o|��� &FI�g�A��RU��!E�R�ĥD���p�ٍ�
��đ�-��{�Ė�Lt�[:��q�j,P��=���������bz���N/|��k�9 ��CP;�?��Җ�n����馗ޔ~�wޗ>}�i��7�\�����BLf���;���_}�;qUp
W}YNӮ����ϼ�`�Ǿ�Ig[1ʷ~�ߗ�{�Q��C;���Ĥk(D�YA�X'�* %c"��31H��%,됍����E�y˦�0r*����M��Z1�^�1[�t���KH!G��e���g\\$c(��8
�'ҧ�~�=�}�A�ӿ�ǈ�ˈ�?!'�+&��D�F>�����ܢ�x�Yy�;�����Y���us�*�:����eZ�3﫣��*�s��It��u����{߄EW�|K1}"1d�]����(�`�ŝg�ft'J �uF�l	t��DԾ˜pgf�G��4�'}�e�;v&'B��R��v,�����KU,lP�qX=��M�^��a"7�!��w܊Z�t(�#��Y�u9��È.�y�3�'>�	���껊��ae1����쨱	m����eh���Az,�KpX�%!�*���H��6� ;1YwN+<%�pnL-���EN}M<�b��*�t�(N^�m�w	z�8�3&�b0��S�α���3�~v�ȇ������Я.䣏=
�����"���������Y��Ŵ�x���Q�
6@XO�3�"xN�k�����~W��+1�G��"�Y����+0wωa�~d~��Z���Cys�B�3�uIi�Ϟ�m�h���jPh��H���m�o9�]M��%�ӏP9�$j�K�֒�)�����r���z���I��q������%>/Z`�k��s��.��T#����r�&�0��]��.�U���R�<v&�F;�\[�J�~Ǎ��q�y��Ǚ?�R�x�m����2�K�����/O'��ڍ�k��+~�G���֬�:-w��+]u9�Jp��;}Ӏ�8ڕZ_��4q�d��lio����&_e���6��FE7�7?�*�zM߭�VeT�*�*�J���g��O>�����t� �V�%Ë�SBA���-XW ���l�~�wFJ�y��2�:� �^!���vwcV�\�#f��|A���4U}S�����ޥ��9)Dj#�!�ٕ���S�=>�D�C
^,dI7�7�lH�}r��C����r�Ԩ1#\8�� 02l�e� LXesӈ	�_�01��b�ˏ�/}���nJ�~���Քv�؝��Mw��wnf�~�E�@T�&��B����t|��8u�H������{�u�R�}���K��2�����[)=�xe�z���#��#�FҖ����%�F,\��Q䕨E��K�Q���A����>��gi��ǖ���J�>|*}�#/6�ܕ��y`�+��������\��I\���C���p�]0V@mi/�m(o�������W]CX�����N�~�S;���mN���[c۴�F����З%v��,��
����u��Z��!��p��o�e��A������H#� (��L�}��#2�t1%m���hNo��|]�Ҫ����U����gUZ��:7���>v�ar�#x#މ�k�lWW!N`A�d׀� n�NDC^�͊��͖���2	�4��`��	kE "��	,69���������t3�4E<.�~O�����u���� ���?�ԅBn����o��16&۶�(_~8�Co2�'p4��\-;v,m�e?��c��`��9T;Ӄ>q֙'&�'�7<?}�#����b�2穀5=~1Q�P w�vs�G��]�a�$2����L�I��NׂtA'y{��22x3|-��w�w����� �A,��Э@�Z	��G1�-z5^N袤KX8/�A�yz��B�Hu߾+�_��'��O%���¾%��m;�~E�r��	��ٗ]p��л��Z=�.�F�k�gI��E��崝;{Fn^��L�[�m�'����WDL�1��k�+'ܪ4(a��R��k����F��T��Z�8�����:A�y�q'N'���f��:�\���H�q\��m��k~i�K�:?֚��%0��O��@���u2�5��sIs��f���J��B�F=X�H[�z�꫟���}�ۈ����ą|���̧�80�+�0�w�:G,����4Ģ�%��y�E���'mt����iWY&p7I��q�w�!񥖋��;�H����k��u�Αq������/�� #�c��4�!�!v��R���>��[^��4Hwu $ý��7������~㳍�U��o�����S�U�l,�9��g�*������J԰�<�g�=𪁜rF���I���[^����?E��=|vH���^�,��,� ��C C�A��iˊ\�C ���^�w��K�.���rT:(p����[[晴�y`a�E�ӇE
�7�A����4ku*�WꮄA�R0Q��)��&GY�qI�9T�s��E�����������������dѿeg~�3�L �1Bt,�����XBW���n�G&�������={�<�dY��>s/�?�����_؛��-ߘ���}�q��ǀ���~w����7�&pgM�;�?�$)��{���"�q�c�v��]q�B�1�=?=��x��N?1C��8��<����oyUz�h3Ֆ��B	X��& �vn�"u��,��`������}Y|�����y�K!;<w�n�Zԏ���s�rbYcw�ܒp9�D����l#VP�A�l����t�n��,yX���bL
��(�[T�:G�F���M�S��xczs�>�xߜ����zc���TiO��\����J�ܡ?�`5U��F�DˍE ��r6���e�ႆ�'v��,J(�}�%��s	�Bp�Ls� �����Y"�r�\(1��
3Q��~��(S��}�,��w9�w�k8�ȃ��?��g	���X8��w>�n�<��AdĕT�S�$��kH�5�i;V�q�7�	:;<`��s������9���Y\���7X��=
"	<Ը[5���7��`�e}��>gb�V�2X`ci�Rc��5�8UePG����D��;���+i��f�N#2Y�ۥ��N1% �K�Ц�"4,l��v��b�W� e]�*uFwc�����&�?�ǚ�l-�n��D=Q!��I[)�EB�exh �k��&�����+^u�i�C-����<:,lR��K0΀�TT��b̰�A���*�]�h	+��� �~��\/ #�REv	$�A9�y�59bA����Z�}�yx(t�^<�\�|�ȼ�5'��E�MG�a�rM���mӱ�=��x���5��D3��FW��!01Ĺ=��鏧W������B<�'j��ޜ�PY/�t��(c��P��ܜŷ�\Y!��̕ ��!V��L�P@�=���a��L]Lw��օ����������>��Խu;��!l���=�PF�te�|:z���;_��<|�<�y|���T�~�E��ۋ���f�x_��x.KsX.��|��꾹�*�z���i����mU��  ���>��l���"�(���QI���a`���?��2'"?P�ȋkK�0��v��� :(�L �v��p��N� �����ؽR�:{Q`�b	w�Ⱦ$S>:2�>{בt�}��M�0�@K�D�f���o@���ġ��e�K���I�2��r(����	p� b2LOq�6�v]��4�Қ��L�+��P��2��|��3��?i��[�ڌ:��GN+m��]�k�5������mݭ��G�[~�]i��^��/�3?�;�W�N�R1y�����a�+!4$p�R>z�|��w�Zz���t��n5�3�������m臩�cs�s� A%���ن��X����_��� ���9���M�H�4��ݙEt6c���ׅ� ��[�F0�G?�^�އq��2����7�|]��o�%-͠ĉ�Ӗ[��?�lx"����Ģc�v� c�A� T�����ȴ�T�����h	Ș��*����jW��.8K�N�6%��>�~�7���u��`P�[�}T^C�Iq4˽�.~��Y�:�����(�I�r��g��ڤ1t$`z:BH�^c�]�$R�J��  @ IDAT��т�E��i�r��'�t9IƆ�gF���o�����T�-���+D��y��+	���J�Kl�1͐�%�
tA�v�}�C0��A0���ர��Ni��?ˎ��. ���>`$����� @��=������#!~���ޜN;�K�%T}Љi��\�LM����l��@�Ȉ�.�V���`��B�%"��S4~$���ek����;�NG�"�!���#t8�5�H�s��P�	�oG�L�3t:YL�
���͉1��9��=N�po�U̡gع�X��:��.�!��{���p	Q���Pw]p�p���$M�?G��aܺ<�.ٻ���7~k����r��,�l�#��ԋ��y����cՙ&&�L���|&q��fYWq�/�n�ݨ�^������c~���45:�1>D%vt M�1�s�3�YO������Fz��iB�5�A���u|C@�i�.�C�4�	?�?��InK�Y3�a���9{4�-9�����:`C�D��+ٍ��/}�6T�{o��'��>�3���/I۶�y��&�U�|���A��CnZBlgm�cĻ��BL�4H"I8�-F��%��A���t����������ok�~(�9����,��ȃ�p��^R�$��E���ZPC�8J�8}�W�-ݭ-+3�gK�%�l���i������*��\�U��*�����W�l�������sUv��	�ԧ�>��k� ��h�Nwץ��J�"9aFf��= ��5t	��\���9�J!
ȥ\���x�ǈݸ��|��}_h~iZ��Q(U�P)0[�M�N[w�N_��^^8!Qd���2��1EB��d� -�ďŤaΘ�q��nP�;E�O 8>�X�Μ)Ճ��-�A̃�u��ӧ���4/� a�x�H��U���������a���^Q��;�k�����O�`>�Q"k�#����d����;v��Ǐ�7���������겴gKN���������y���fC������v�=���>�9tm��/���lV�!M�F��D����<ֶKpvV�k��^������w���W;�1��CP�@hƤaQd�;��Rwj]l������t�c��M0��t��	B,��׿�D�,����w�{�;O����TF"p�h��q0&q��'c�e��� @ǒ�T��*�m΁$���RE!�qq4K$Lz��r��+�ee6�_#W��+^z���;���O_E#h��/X:X�����c3�`uS���r���%�=��������c	~J|C$@�0<B�&1�(�`�
�H��{�ܨ�[77I�R�e�L��F}����߈�F�����-SX�RQ��Yk���"	-sg�O}�!��?�FTZ��~��=�b�q@9��*���u�����2��D�m�45���^	2ǵ�	6��O+��jX�m�Ӆ2N��Ǎ�u��(�M�,1�P���:ႣX[S�y�:v�y~z.�"yb�)n�W��P�ؐ�S������������04�˘�WD5�Q�ׄ�BG�'N���q����O�~=��B �;��ݻ��k�?��x���p��.��Y�c_�:������mK��y��GSO��<yb��M���8%6�zI�8����K��@�?��?�]]���p��j��E�&[k���I5���S�8�JB��_'���u��R�K����SW�N�RG��2�F	�勑f���b�X;:�CV.5P�J��7�����fpu�XE�5����a�wx`ܹg����K<)1�sҹ�>�c�V�v~8't"������я~�x��pZL�U�w��x��59�*x+�Xb-Xe�_v3�R�ɣ��u���}�w�_˘�n�Pt ���%�Tv�W���?U~��F��+�.�oN��NU~s����y����<�j~��v;��ط\��T�<�S�f��=L�9�F�11W܆��>8 ��U����$&q:uXT��
T세�!��=�<�x4�@��/
�q�x�ecN��4��LUO}�9��������֪9�,��E�p`uW�5hlj��$��*h���H�I�ʨ���>���ه�WKO���1��䞶��0t8���������G�]{�ϣ��Wn�?��I��e����$�c����Mצ��O�-�+0��+*��� *�X��u�u���{�B���S�����~���=��굙��(:@Ã=E�j�f^дǦ�	E2��=����z~`���q��NS>֙�g���q�C<�G9EД�yh8@�J*��q�U ���8�HB�}p-�"�_�:%�C9�,`
m�<�|�����h��[�Y̷�x }�����`��J��0^�M]�0Y�:����|
��o{qz2�c�Ǳ�c���^�o���-�p�|�HcU���4f?w�=��Z�#���tt�a[	N�x[T}�}P��"�����8��OY%e �T�z?U����T��\����x(Ǣ<�j2Ti�dy���m܆�q�*풶�+$�H�s�WbϞK����fLzSa{x�?�_=�k�$�#3�Y�BI��\+2�HC���B��&��K����a�0��&���-"����#��<Xrņ�`4�g"w�%~�+^X��4��gэA% "��~�!hk�8���J΢C��UDΈ������� ��S�JDq�t�8����ӧ�0zw�e �̛>mg׼Rrt��#���(����� ��9�����UT��6,�{ڋ9v�lZ�����EL
Ul���V��	m�Ի:�X��hg�؍���U�[+���Y](Z�=ֲw�W_�^���.��c�1����'��� ��2�}��Ky��q�sn������ȅ�����o���D�O�pH�
e�!h\���(��^@�7Y��>z��$6�yH@(��"}'<�M���;RpMKKG^n���`�j�7?���c�F��O6;;%��,Fz ��J��92tT2a#��ȶѷT�a�|����2��F�"ܓ�lˬ_�w�j�2�WV�
�9�Y���h�cr�(�9�8j���J��\�V�h�G{)f�hH"<g�e �������	]FLy�_�����p��c�C���]��I��(��P��
ႂ9�}5� B41W#ZC122R��0_�y4c�	-S,A���G����|�m���y����[oE$K��D��"1;z��	�Z��;�eTCʨ�����ܔ�<<P�w�C������9�<诨��2��t�7�s��s�|�3�}nz�*�z�:�W�W�5�7�����g�wL���#�v!�e~[K���`%�Tm�R���L�{0��}8��/I�(��� P�6�9�{&����H>n��E?�'�X�H�,���!�~)(0u8�=4ӕʧ��I:�Dhx�̓u4�{���Ƥ�< �#�����c0�mA.p��DF�?&=ec3gf����,鰶Y������%A�`{/����8�KS�c�N����-m+DK���z9"ʄ�Y]Za�!�`�^}�R\�C�Ό��nw�%`�d�*.�[0�6�Xu���t���"r ;��cdcUb����b�C�l�ױ2���;S��l�.d��S f}�������w�֧7E+�Z��hӁ({ޡS�q��1	mcǊ�J�.�G;>reֵ"R��?{_zë���w�M�e/�#}���{a$@@�剴m� ;��b����/}�{8u�ҟ����wav����+3(���ۂ��)����T�W`����^��+ ������^�Z���O&�R��26��y4��ϛ�6_�vu��\��T�z��*u����)�m��m���s��4���e[K�#w���YB!�Ѵ�1�|&�T��ro��P�V_��y�� �".���u3���� ��c}\ �K���],��$1�N�:H�)��3op����Y'�ʀ�P!���#"���1�}�]�n<��_�;k�G�ē��b�c�=������\���;Zv�F5�5H%�&�@����ʣ������y���{�3�!�`��f��Ї�:RKP��Tt�}�B�k�	��;�:q���)��u#�(x�aw�U�$�EC��uk�F�ސ)�"pt�Bg���(����N � � �G��O�d����5�O�oiz�9~!b^�tq�����X̒1���9�l1���T�x<
�\�+W�	��6g��S#������o�EB��IkI�pg�!B�="��wj/CY�~�nx�R�_�/�+���Y%m>%�I�U;�)R�[ݦ�K�LP�1��B(�n�X/�� ��nR���:fm���'��taL�	��|�	�����ܶ=,;��r`q���!�S��8|,)fs.�=��-��d0z�!S���:�Wu�&'ǋ?��?�*����J/~ſc>u��YF�A�����c⎲�H���U����^}x��'���Dtiu�7<6ޗ W�o|V�Q��Y��:��T���J��UY�����߫�V�V")�h�l����w��cW�5��� �rG�|��?�w,�v��Y~��D�:C��U.H�h��|�:�'�Ǚ;�y���^��KS�'Ve����x�����a�R��3�셑���}Q��򝰱)`���!p1AP�`�ǘ7B~�.c|��*��XTÄdZr�"B�%�#��j5=�n�Ɣs�bk��R�&&Ɏ�����V���9�ュޱ�9+Q�:�	Bj.z�v���b+v����+�K���w?����i�K��X�NH8{2|�'kw�T�����������`����i�11.�G�I`'�0����@�X��U�P �6�xr*�:� ������EjL p�1��K��X�>d\^,�C���.�;�r�����4N��x����wmKkӟ�CD70�� 
�������������Н��S>=>���u����O���ڋ�1��'6�  v���laj�Bc���-��b�@�����d*�����7؈��w���^�ҫ����1��W����FZ	�Bb<)W�H��°����9R��1�^�K$��E���꨸0��2����b��[A�hm��ď��m��ǚ'[~||G��!ڲo�.�#%�#'�2+.������$�-�f��'`O�!.D�5�}!�(V���N`ΚzQ(���wr�p}��"�!
�*�.@���Qv)�s�^X�Į҉�������s��EL�%��7�(�%�A��)!��/��w9�H�Dї@�z[�A���Mg;F腰�kH�+��=��!!���(��GuX���r���G8$�x�ȁ��\}���IS%hoJ��y�,�d�S��e��0��M�`\�ݫp�al�_	фC7�,
'��o:"`Ł�Y5L��Ի������r����: Mw�v��j�=� I
�Ҡs��\���*U4]�L�܄C�m�4�hp�]�Ք�����$�2�Q,޿���кCc#iu��"f8���d&�,�����$v��E>�4�c�`�V0i!ƣ,F�D�N"e�I�i��)�l<�0�{��H^tD\ ���i�G�,����& <�m���=ŉ��J����j�@���L����r�X��G��[�b7Հ��p���nX.��Uځ�c����9?��^������a\��P5s	t��Jĳ����z�K�ߝ>�wo~�����>:=VG}���8�6�<��M�'u�7����1Gs�F9~g=�)��/��` q�bb	c����$�+��Zwߦ4����m�r��!03��o1���bf��v�E7�s���N�u�r9w��1���!ș1�>��`���X�RV��4M����Y���<z�L�An�s<�.&�����H횎��=M%�f>��Y�y���H�I� z
��p�t��.��}�X�>v$�M�R�%LqZ�4��͉|��Ø���{�[i�S�N�?0�SȔ6C�-��J��E4� ������]K����❖Կc_�<��)E�?Q��:�^��}�������2�q�4�B���|n�,b�F�!�ls�n�im.;3QF�	���(b��-Ȓ��EDU8��63d�T+ϙ�H�1�D�pE��ܨ$���s6H�4�2�� ����G�s�I���Gu*}׷kz�3��~�y�}�>T��t�r�����ʍ���l('�����_[Y��ϦR��k���)��o[W�O�虳'Sצ��ӏGf�!��p� 94�vk�`G�]0v��t�S͉�^tb�7g�W��չ�y5��ZT����4����ߐ�(Ǎ� ^Ze*�����2�s9E'޳�W��hAd�0�Bu6"e�V�YbB="�j*���1�d����?�Hr��� ��6��� Z�;vd9<��IX�M��uU���2Ls��Y@$��hY��܂�����<�.O�	<7���Op�B�պў ��L͌��%wЎu=+�)� N3&�&��0N��X�5ݤ�.��ws�5D)��V��E�/B����֍�9�E`}���K��)�D:!��$XY��������8���c�f�,�Ւ�, 6�b�2`&���iε^8O+]@
(�;�I2&P�n��^���4QO��6G;������Fgr���J�uS"�,���H�/C�9^��˚@��!N�".�p��m ΉR/!Sz��S*QJ/�b<E״��>��Y��%"�]�@���?rt��3)<GDr��g���b[,^Ћ������3�ڱT,�"]�����5���ڻ�Q��#���
>F�&<�¹�d���Kg��F���ˇ��1�F/����;���.G(�n۲�(k�۾�ۀ��(A���Gοy_Ğ�n�zL>Cl���?�۷��,�&HN�U�u��冃6����#�7͊+Y��9hin0��	�Ҏ�y'�ݴ�X����P%d[����إ��8�~�2�c���G����(�|>��W�W�չ��+�w�o�����o� /tև`��%��3�?%�Ov��!��p�d���%Rt�ˌ�0 ��^��A�<���bDGE�����ۈ@�-O���j�芲j��7��h�A$y�&�V<����N~�7� �'���RJ��٬>�^�0��
���L��k_zC�f߮��.��N�+_����c��|<�u h��1�;&�x���׿�E,�Uv���&X.&��	�������o����Wݜ�x�=����i����A(���]�����ǡ$�F��!H��y2��/�7�mw��w�}���k-ܝ,��f��Ǿ���w�J��߆ub�9�	���ހ�Fp��š�c"G��+]�(4��iDO�1��-a�PF4h����s��á�]���6ܞ�ݿY�֯���=���ߞ�����8O�
��=���o�
�0�H1����p��m�����M���e��Ϲ���g"��0�By=��ܑ��ƯK��;���$l1��r�g���O�xM����WG9H%a�Έ�`�}�4�3����{�4G��s��YX4{��k�'}�L��S�S���%�W�%F��ri���5�r��hX�3�SꗄFe�$�J��~G]bȶx�Y�,�!�#a!��}��uD"bE�SD&�����G�CYDm>�Ur���DQ�27�q�E�;�>\Eh]�70a�qu���d>E{���P*�K�)�YD�Mݦ��;�oZ����Z�A��.8,��J?�<كI��%�B��Õ���b�JR��u�E_C��6Wa�Lt�T"sm�'gt�:���L�R|Ja�-ל
� ���%�[�@�_��%Z��L՘�Z����z��nt)���]bo/i�ߧ?j��ao���Jc��By��l��P � R2��B�`�;-�#ǄrR�o5�B�
M��S4_��}��t��#��w�!���.�i���D�cM���8ZK��qG���^߾{��A$b|�x�,���Kr�U��}�ܝ.�-Џ��b��v��E�j�M0����2� 8R]��5,�b��V��
��&�N��-��:n�sO�����:��E��C1g�4�@�	�d�(!�0�SP|iAJ�����9��eL��ڑ#G�n���v�%y����Q~�I���ŇU�\ט��L�-�S>�{-��oLC���c�X8�d�r�p����|��P8OTN�s!�Gq��9'��S?��s���x����3+�,��F:�9l��Q�Ug�G�*C��}�u��9���W��\�5��:�2������|`
2�nH���l�VлY"�b��	v�l˭���4�l����)����+F�9�H$�ZN���P+�-�i��_��o�<y"ED�?LMI%���r!X��W\�U�⠑������h'�A���"&TPYQ5�\�_�t)��#d2��;�uuvl��'N�������Ʒ갈�2�m�+��������1��q���=�H�pFL1�{m�j(l����H�͖���}`���/ٙ&/L����|�U�ԿA���?sۉ�����H����斎c�x�޻%|����C,~�=�M���D����'�s��v6!E j�B� 5�t�;ۍ���g����O	�(��sS!b^�{(��WnF�y0�DP���|9��{?���}'�cx�&�۾��1O�����L4�(�g�ώ����O���{�^��8�7���|oڂq�&��W��Q�FD3���o�������������[�?�CE�}�~�RzQd{lu�M��lQ���l|u�9��? y���[�_�gB�h�ހ�'�zf����=M�JR+;�/gE'��K@`���K��E�<�{`�]�iA`�t�.��9�A������x��H���⨨/ʕhRt���-�������7�i]����!�B,�U�V>,"�}˔H�����}Z^�?�X����C�W�v��3x�#��7S�Szu���p�`i"?G߰���낤�G��4@�D;����APJ��Eh�+xF�%<C�b�.ƃ5�g�/ؘ��R'��[�y.co���@���|B �m	ج�Q�^)I��=D�R�ؼ�I�{�c��\%Oy���S¼FGOsr�Ɔ��h�޼�<�h7<����A	�o�j���Z7Z�R�����8Nj��ZǼ�H����ߣ���3RU�Z�����U��w�};t�@��)Do��?�����g\����	D|�;��w��p�/��-��*\LO�+H���?�.�qt@���TG���QiewF�x��P�ς��F��¾�8���~vw	Dp����[��l]�rk@�J6����� X�S�`EΏ��t��Ӊ��b��p�3�y��ĉ��=	�a�t~��)`^A��oz뎍
1�_,��_����?�3u����~����7���P�[w���<>��Y��4�ߥ���a�݆1�v⻝?��dn�U��N�~�l�s9�js���s��9���t﫣*�����孞Uy7�����yݜ�}uT�{�ukWK���K�20�y.�
�6��1#\Y[�i z���u��'�ko ���z퉲�bJ;�T��I�����̎�|�#�Yj�&��-p�(�A�B���%"w/@��cڄE3�D�>O��GWE�?p�:%�_tjSw�K���|=SO�9,`�>��ϒ��^�De��ߑY���� !8/�^Xs-�����?�_r�X�������~�s��x��B\��>{'�W�9�\:�����4[L���}��r׾�i�δ��.�*��>7���ڶ�Ý�5W�C�N]������x����y$Z f$�;1���Q��?��'A�[��Ư:G*��E������0l(�t �/����W���b�ݖ��W%,~���1���ņ9_����K��s"����j�r�Ui�Ś�q�*� ݙqqP�4�ۊ�9������&e��8pp_��]��7���)ReG����lc[�e��"�m�pD�I��p\�	��;���;�w��XL��i�o���w�>�J����W(���bq�:�r~����YT&'F#l����Q�Y������c�n,"EI��鑸�0
�0�� �n%8)VpNj�W��w�t%.����H(��svGk��O�D�7��}p�\4\���e[7Eu��"��<�9�9ۮ+>����ǏgObb�Btt�K\���Mi�d��A�)��ͻw�	Fvf�<D��S�R�[8�D}��:���C���u�t�7@��L�g�e7Db^����s:R�2�E���M�y����	�-pE�[�!M m�	�.�jb����8|&.�d��� ش��8 �����DHT^8�P�@bH�:��&r��Pq����D~�x��4��V����7"����37j��jlH�f�5�=T��:�@�Ϸ���p�rðC�S�����$nLfӴ�oo[޴ykpXPԦ���c����E�����-��,���֭�����B?����O�G�ħ��U�9/��p�C7Y7���j%��Q��;��{2�U��C<�Š�G��K�����e1��|�w�.�{��'�h#�p�R��B�.@��v��i��E迹�����Ç�G��P!}b~�I�xzjj"��y��I�n۶=�FOL�lҭAt�D7�ıcI��8q�`���cǎ��s���z��3��!�Ek ���sU�M.R/s��VQd+�Ď�� ���(=�Q=n���t��<�WelL���=k~^����>�>�f[3UJ��`���@1D��6��� ��\p�d���ɲ���>n�YV�Te�ڔF��d&
{f0�DL�2w4�K�_fQ���]KpA��ԚI�%Ri���%I(X5��:@$�6�Y#�S3��T~7'�˱dR�;މ��7`/SL���w�����'nՙVZ�7� ⁅�Y0�Av��%-I$�����\��P�6~�	��҇>���%/������|�y���?>t_��������K����Jǰ��_�l��k���'��t����=�����}mV�by�V:E�+k ��r:62�>��O�#��b���k��~�w�@<��a\��P[�K��@�ƽ�O�[:�%���ȳ�P-{Bm�t��N��~�O�gQ�<���~&}��_L��{
�Na"=��"�t��83���S��Uץq�_uv����Kh�l���y�0��:��J��	>.���Q�3�8$�ɗx����Ϛ�-�Xv;ހ)G���Q�'����}#y�Y��:�9M��#Y8|,��Y�}����~���ޮ_���y�mwq��JQ�����[�Ңu�J�Do9�@G5%`��w�8'a���w�*��C��s�籰;�>v���`y|#�eH��b�sF���-r�*��b�#����Mn+޽{7.N	s����ɨ[��.��^��TV�@������!�cl�B�D�ŕ��@OH#G�EPg���� ;l�8��������HD+�5��ǂ"�b��E�	pe�7mf��e�i���L&Qk��|�֔�bs�!!��{�����M�5�IP�aI*3@,)/�yi���E�tll�p�|e��bJ�`;�1�t-��x���d���Ÿ�������C���2��SOH�1��9�HM�}��K ��e�r�`���E�l8���b��^�����|������{�M����-���g��K�k�փ�}�O'߇XA/L�6�!.���TL3s���������D�	�O�0�c̏�%��r����˜�TU.���͵�����8ė�X�m���ثȏ��Q�.��@n����߰P؞�8_,�q�]���E`�1���C�z1����k�����q�ãX:68T0�'*6̹�`|�����ΟJ���?���EG�S_L�-���-F`߃�r����bW�0B���\dó�{ę��� ��?N�(5��ӿZ>�]|���]����K�y��s��ſ��U9��W9�*��~����V�G;�}�?d��ND� 4t���2Q�w��l�(����9D`��ȲQ����tfч��*;�� �"���4-/��d*;�-h ���](��`�BY�����hă�/�|���?mcDQ�	.�肜qZc'��ޘwa7:
z�]�hֈخxN�G�E͆�����@�8��~D����,��[������Ȣs�����XZ^x�(�{S+H�� ��S����K��?�bFAX�-��;x#^u�qD�K���CX��b&\��O���i�������0��}�Vk��~rԓ �BG���
��ޢol %���~�{K1�EN�}�
e7;�E�.������0%���V���y(��rn򅀥�z�����)��kxF�"n
�3i�NWG�Fɰ�i%\,�1�ky	0���hP�l�1���ZI�+dX��#�������(��*�:[�cK>.ig�T����I�ʍkऺoz��$>�T���~�A���}��Q'�����M�vw���8Ǎ�h:W7�<1-��ݥ�Vi��Zr�\\��9�����;����J4�D*�GB�t�I�>�@�PQ`ǲ�Dl]-Ϻh"-A�x�ݴ�I��"8��	��+�˰>^�mE[���43[<���M
1\���gOE��C�LNIx�o'F��:���
7�6��+��Ehse��X��B
ct�X_��6Dp>���c�V��	$Fm��!AQ�.�F�){BV(s�W�63��q�;��"[��; �7ii��=�]6�K�s�qԈ�kfSeEc�)1b� l~]W���
`c�K��P�P�pm��c���������~z�7������7p�1����X7p0K�F)�g?$&A�DA�@��7E;"�yj$�#6a5'n�m7��� =vL?V��xun����`�?�8���E�ݮ�o�s B���⢖%8^���X����&jiNeW>K� ��',�8A}�;������y�p䋯"!�n a�h�u�w~���R]�z�:8qv($)}]�D��I"I\�<`�>F�
�\�aI#|Oܫ:������y縸Q1����9"ד��a��g{b#��֮];c���*c	q�V����Ŝ�{��� 5\��_w]9�:G!49:�ws8C�xV<��H�o��&�І5G�
�g����cc��{�
�Uzu6�k�U�f�����W��g^oL�xo����D�bnn�R��$^�&�>��6���%��D�q��Һ��y��,��1Y�l�����������Xנ�ټ�Y��P���,F���X��ؘ���\�:Ay`�1g�'3�����n�+{Р�n�{,��d`��,�XQ3:Lʆ��>P;�.��@F�x��� �3K(�5����X[��k5�� /���s:�H۵�����Z�!bDL ��#��UW.�:&�"	Z�2&�3��e����Z��Ch�W]dF�����e%jig��_C�~� ,f �a���-U�`s��$V�-�h������� uԨ�EVBS�@����Zݒ��YB.�m�<{4Ζ�s&| z4�E�F�R���1�a!G���s&�E�ߦ�䪭�;`�����^��n�S��ޟ�����%\���[��7AQ{+M��z�5q�����F���R���H)ߨ�6���Uz��SYj��9O󵙟._��ʿ���Iq�l?H ��?�����%j!�E����A�r���a�"d#�Kw�|.{L�n��;�|��N���N� 	���;�^�o�qD�"<���a�~O��9�/��h
B�����*_�� zF(����,Z �#ޙ��(H0T�BA$Ewn��4X-y���IN-��������<b��y�ޝɘt��$�Z�DD��&��%���d��#`X�C�`p��lxr� �pO�	��0�X���,�@�Q�e޲
!��7�&(����mH���.D!�����{v/�)t�p@g�@�,6��(*��5�?�K�������op����M�'�NaJ�p[�j��,�9�&D��/l�9_��q�汦�����[�ԍL�����e�&|YM���aj� �ݶ�$-YEf�f|߅�<x'�wgGO�k�ui:��O"�?���c?�n|�Ş��1@���ą��w�J��mw���/#|˹t�ŏ��A�]�/���c��\ڼ㒴��'mꇠ&�� ��l�,f�?�5C�A뵸���bֿP� � ��q�!�Um��6ݑ���?��EXG��H�S6!��e$��|
�~��n�Hᒽ��-��VL��N�_������|�3i��-!V�766V�~��)cS���!�Lg��Ģ���=ᴲ��6�pa�M����P���5z��[h�8�y�2�F�˭[�.�>� �LĿ��s��X�}}czsލ���������N��n�F�s��B�\��&{���45�&~SK��]���γ�s�Z2AB!�lg}��H� 8p�Dw�Eg��)����D�@h޷i*�@T�����<'˕�����SwTR:99��S^�M0�_ͳL�����ͷ]q ���!��̥��o-�;\�|�� r����gz4���N/�������3Sx��C��5L4vNp�0`[_7	Ǒ�])�cq�_h"�W�Y�_-+�3�;V��*-s���v� O&�Ut��{I�8�� E!���p�4.�zD�#�4_��d�ri��E����g7P#ˍ޸�����l�U�U�*�bJ�/6A��)y�7\��gcpr��(U���`I��qݯ~1V/P���g|�´� ,���S4؊�	`=9�U���,�GB���1�|$;/��}B/	���4��~T�2!�snN�2ViչJ���ݘ����U���>���*o#�Ԏie��1t\M��#��(}M'�޽3Ϗ>A�"ƊL��3G�mJ4��+���nN Ua7m2�����V$l�+��2tx�9o=�����.\2�%��t�*��$���� �|%�p�+� �r���B�'�Wcv�:�#�-^���ݹ��Ⱥyx��?����4oV�@16oټ)y����%?��0̈́��	HZ�8����؍�	G��A�͚g�R)rCV��y�8pM;)Sp��'r���ί��!#Cx���-P6�1�)_Q1���x	��e���l�Ե	�<� �z�S����CA��h�D��������M�����.�_}�Y�	����L ���Ï�W"��ló:_�Hg�%ƛ��3�9�hrpS��zS7�#��!0�\KgO�f�Yԇ�FE�T���`C�PL�`?:rj+Zӡ<���]����Y�-қ~���۾������Γ��=�X2�0�������{�Ϥ{��x�u��O��Oc��z��ٚ���,��@�3����γV�0���#��+�ǿ3��S��Ǻ�<��szDg��n����J���P	kC�-M��@Ĺ��Ic��y���� ���Bvo�S*����}�-�m�m����M�V`�� �_O�gN�^�<��O���spq�ݗ��e��-��3���8c���zP�l,��*�����v*Έ���A��N�ն���t�2��cn���\!������p�uuoZ�us�*�:�L
;�[S�eٖ�TGs��u�;���s˩ҫs�}6D5�<�ڎ��1\ߡ@�̰d���gT1,�UDQuL�quТg�:]������Px��C��Ð�c��J�My࠹d����@�V�����b���p���9t�C3M�I.��m��ҹT�1'� 0,�%���}4���~������38I��:����@q���/���⧿��ཤt�ߞ��{� ?~�N�+ �.�� 9I��P��pJG��j�&�z�� K�k>�
�ֶ�H}�;��|X��4X���$(|��� x@!��*s�㴌��#��~sr����">1�������s��R.�
7>�� ��>ވ��ܥx  @ IDAT�+ϼGE���%s��L~��QE����R7ax��0� ]W�Q�v_�p��W�S�t�C� �W�%�3,�j�Z&gݿ�߶FVEr��S�������z��8l��O��*�z^��r�﫼�O��J��Q��s� � @⿻Z�l����0"p���Sl��ҳ6DG`4ދﻠ��/8w���9`�����4�]/׊x��Mpg�%�2(3��LyAXI�Ͳ�|'�/��&�[�k^��3��v�:�ft �\���]��Ʊ���/?��&O`���^��V�;vl�]Z�o
��(������1�?}�h��F��2�\�p�� ���*�\��)���Â���ۘ�r�! }�L�[I��V8_]��e�L�SC=]�k��#�"v�-�HM��u�[窬���p{���Y��b)��U�H�3�n����Nu#���p���#�?Φ��v-�"�������r�p%�X%e��%rꛯ�m�7H	f��1� *���H�Gł�����s��z�3Q������
���|���*!�������"IDI�͛�q,��ڞ^����X����?�_�I{����`�嵯�8K����]�~�G�}M�	����I���]yi�B1����c�.�A��������I���i�7 ���O$����(��
�"�.���)�f�u��YW�].�����.�-L��ݓCߎw��O�:Ai����Mߍ��up7��;�6�'��;�#��Ip�������]W\q�广O�Xj.,��.=��}����t��1�S4 ���0��.�/P}��8D����J�(Y�&�~u���[��pm��w� ,����{�Í��35.���N�=Y������O��<ݳ��ah�c�f!�Z�yj�_=����M�\_�.v�+��P��^�
ja�i��p/�r�k*�a�6�.P/��ť�]���������� ��%T�"���tQ�nPd�oj�A;�rbo�4���B�`°���/�'"1���X�Y��"� `M=ID
B����
��8x�$�v�L�2\E�x���ֿ��DX�[�Z�1@�5?&sC'��`�:�ESu~&DL��9X��3"p�R�(Fkm�h �bg,�P�
,LM�C��7��a��<$��	"�;=���%�DL�.I�?��G��~e�x�1-hN�>�"d3�e�`-_��Xɨ0u�*�#��0[���wQ_f�*��)	,�&%�`{C��9�#��P�m��bp�ee�5�-��%pa'�ͭ�O��S�Iz�Q��>l�n�\�ٜV]W�T�*�suk�8�����M�)CG�((!����"�y5�~�S'1��ցG���o�)%���+bD��y켓�� ��(�:��b',iv��Y.^����H@	�[T:JV�EN��g���@Ã8��ջ�	����3K�����&梞�g1&�!���'�Ĕ��,��T������$��y�%{C?�%/~I>{v�)k12C�+G ��WA�wl������I�߿	�a]�Q �7Gd�I�����p��ʩ������&kL�0vO�X��r��&�� hkE�po6El*������p4�OxjF�����ɢ�����Ŭ����T���>��{^���@|@?pC�H��"��S1��xx�mc4« �1RGk^U�Sx&Qn�pDԒE�(Rҍa�( �J���k��b~b2w����E���C���&O��*ctC;�%��a�^K� �V�Hޏ�� �����~�gޛ������<+�-��y�ϥ�N�O���oH���+Z{�����\��Kɉ�[	:��;��1���#`	1��}����'� �p���k` 3,=�R��'���~7�������/eP畹�y Q㡃����)� B+���5S}]��V=�ѹ�p�*G���}��S�o!og3 �(�ys�����` ,*���{^ھu��e�	<����˚8W�S	1���
����7]}p/`��ɫ��&d�<��,�0���[s�ss/j]��[^�?�sg��4���c���.ȿ�!2�z�w�kӫ2��i��\�7�c�G���{�_����ߴ^�3@"HȞ�x6I�Y˶v:���Pier4�卯��8�=ujQb�E՝Ԫp�{ E�$Z�=ilh���;�����R�7��e]�d4�*v&�ó�<�g_�@�Y9���� h�ϵ�<��/!����e�,b�N���6��R �~T$p�`�F�^����Ik���^�}�(�(�kc�c�(GB�/��#�2t�N���p�c��̊��*GM��jml�����iQ �#]J%pV.:�	�`���"�^A~F�g�R�'�HY��A��l$S������2��9ѡ¢�Z�����;�k�BM�
>÷K��W�%2[U�O�n)Z�!@Q��`�2Q�g��-���ی�(B�E[�<|X9ED.@q�G����&���f	V�	�]�@(���9o��S�g��|V}�w���*�������l\�$�qW��yH[�Ic/��M6�mXΜ:ɣ��%z� P�3�ݟ�8!�np�L'-����{�|+bH%[�I*��}t�j��8b����������#���ߗ�h��� ���b�p��:T�4��Y0t������K &�
�mř'��'N>���Bc�t�UWŦkNE|���Bɘ�&�9E;00�?�����i�=�бkCβ~�ˢ	�pi}ۇ�h�E5�wx��S%A��1�-�ǥ8C���ş�<F_+�$u֠0=HHD����3'�X�v�a���}Ǟ4>9	� �ا��	q��&P���� �n���FB���9&����1p�q�6����R�F�R�M]B���L{��C��ܪ�u�B-p8q��o�����y��e��JtC�)F���K����b��	��5F�`��ϪP���}l��'��'��2~2�7m����@�sSO��g0��?�P��#G���r޵�Pqϑ������?��o+ڑ���<p$���
'�Seh_�NFY�� ����ą��)ty�$���6D?Q9�>ڏ�<:�`�g�[��E��E0����q�<�SG�֎sT�Ʊz@H;:Yo�|H@��fg4�G3~u��a��Vg��=r��;.���4v�\���s�x������m�fV�M���=pO��ګR'�#tlRO/�EʜK[6�ϥ$!r�<����ȏ�<�D�o�)*jz�*q�&�D���-��:���k,6�l,�_t4�k��e>)�ӫ<�s-^nN���oma�,��ۇqyT:�cN�A�?Oġ;��4:r&��k��=��1�4b�M��nT��%�U��U�9�K�y,�{v�<2�<-!1��E�N^{�\��fl� 5z�䰐NR��3[�3)Ld���A}�@w`5�n��P�yτ
�%�2b����U`�ΖN(��Ib�Dٵ�p. �,k��
X�)�jԩ؊0���,�� l� ~q�v�[���Q�;hT�{P(o�V#� ��@�W��yY���c7����L�	�ƛY	w���*�t=���Q->�D�#��to��%��};�*S��0E�H��|�%9R�}䊑"A+�)�+�,)6�"-���h+j㼪��������/��(���nhB��Vdo1|U����Yn �� �xY醠G��@��%q�k�����x{pͮ�0w����fΙ3�LSB�$d��I�`c��Il�8vn����'y���<7�88��$���0`�H4	�I#iF����{��}������H¾u��g����[��*a���T��mӳ��e��lU-�P������=�dj�W_�˫.M�=�#�󏎌S̲+n<J���͙��5����-�����4��9/�?����N\�;ޕ�P��oa�*�:l�ʵk�p�W0�[�|3.y�IY���薇Q�Z�}��S���!N���U���6�F�^����lh\��)XGݿ�Rqs�>�3�p��T8�;�|�a<��g7�'��9("t�'��[��z��@ެm6d����`�aP�*fb�6u���hE�utu�S�����zWgge߮��6:�vى�I��Y�p&�� �hi�%; �677�uBmڳ{G~�����sW�M7�,M#$>����.hl]��NW'@�P��nO�'C*�,�"�A����$C���!BL�2PN����8fM1��IPF^�#	F�X�1����.�B9�V��Nw֛�*�'�v�?03� ���0��^x�&�}��"���}�����|Zڐ�Օl�A�͜�1�F?��Jx��8��8�FSP�`y����2��[;�W�W�*sT}-כ��ۓ<��I�.�C�q�*2�4�����\�s�\;&H�fS��=�P����α�1/Z�N�a��h9O�vx�d�@�ȑ�ln�3��Mjh��"C������׆�^Xn��I���Aa��$4�
�l�fԼ�l@��Q�:�t���;�7��M�o[gV`{sg�n��s��&D؏?�d�Xyi��lN1���C�l\�w���LΧg�\H0GӉ2�u�~3sSi����7����k��:����WY�K��%��,p�,m�Mݗyou��E޹���H�@{�P��;q��4T�k�UE�S�N-�;���� ��9X���9-���e�l)����6-y��fV6?��N�M5���k�z���roF7�P'�E@�_װ��RO�C9GH����<K)����F�ъ� �`�.eox��	�0J��K$ u!�@�`�qw�gAB�e��s֖�]�|�s����Ú�\�������|W�-�b�#�����%����-	:��X�=���"��X�mh��}��|l9�N:W��X,�� ����!���QdC��]'**�p�hEnsv@U���I+�j�) ��짥r�yw	r�?q�(%XbK�/'N*�� �Н�\�-�$ �:�-�w�� S1���0�xW�P��cQ�AR��R�����ŰN�ղ�6QQGǧ❧�z�BF���� ��@�%�K�I4�M�ضI��5iiIP�Ħ(���Ug�v�%
��|DL�(D2�M�Nra<�8�
�Ȕ���\r��nn�D�6�6z>D]lxA!3��'��x����8��e��[�O`y/���Z��i�V�\ƭ�חY�\Ʊh�Gv2��o^,t�;�v��vߙN�xV�N .egd�y1�"��M��3��&U ��Q����~868�F��"��S�D�!��������,"*���9�mݭ�?��b��.(?���$��fnz��,rG�Û9�������Ɇ �b��kW/�Bh����ھ}(�~tD:��u������?�z�A��Y���j��eډ^�.��!O�$�ZȀc��"�Q!�.�Ҝ���9����*�����c��BL�EH~<s�GF��^yK"N�P��8���{��cȗ%(;��d���v��n�� ����	kM)F��]'�[q�ﲏ�U;�����r��^��+�C�j�ɾ�M((��w\I���T��RW�_ 4D�X-nF�6��BิP�<:�T��*U3���k�/��-7� ȍ�BR���n=��Z\���ܰ�";,�T�� �o�NWG��#7b�ߏ�AN.�](���o2� x���E�Ć��z��mP`�����݇��T.����͍���$ �$�Hʺ�ӻ�pۥFi���a�)��`�um#��7ҧ�k�\��m�#�AFm5�s�+�s��Ce�E߻��g��_H��@��.37�a�-1?��}V�4V9�v����N�\�g�p���͎�8KW`�u{��S���������O�F�7��]M]�X��@�tL�^>|u|��k�z�S�x��,ٟ���o����3�Uq����ar�8"DS�k &����0֎�VG�T�����a��"��q���F{��K��@�D�	_5�H�c�X�2��Y��p�k��D|/�`Qc��5��[,�]#��s�/�A,&�E8]m�Ĵ��_���� �=��h���E��1W������O�,�,
Z�'7�@v�$*�4&:YE�3e���q0�%��;ۡ%Pt��.̧ѬiWQD�S��gτ��-@R�4�قI\�����f�H�fY>؄�B� �=�v��xb]S���̔v�A~����+ �6�V���N,i��bH�� ��� 
��e��)�'�IЏ�<LcT1�)a�;o`�Ed-_k����Ⱦ�>�f����d�<a#��V���	-�I�'� ��ƍ��iLC(b�Z��Y1j�ʷ��͐T�Z�9.q	���CV+�;�[�\��5*.�A Ya E�O�"����KĈ�����l��f}3lc�Lc.12��`s��D<�� ZʆX�s�h����x�;�����7"�iiP�d��u�;�"������3oQ�i����P���lݵ��q���PW�j��d#���K-�tsH� ��=���v�2/� �e+c�F�090F�me�m����Ѩ����勁�<�W�f�>@H������>��29y]��PD��/��/��B�ھs��(8vr�Au��U�W�F�5t��G����0�%������
�>(<b�ug	��K� �����%�V҅S�9��4�ᡷ�r�R疦��h�����Hߚύ�gǎ>%�'{���yX�O@e�^R��b�R;L��|{w�����ҁ��ӧmK���~��a�I��x�,�Ç�@����~�m{6�����?�t6������7�&��{�7�l�m��w�G'�}r}���L_��{i��|63~%���c��؜���Vh#�,�-jxW����"Jo;n���#��A�1��Ұ���ܐ�4�i +\� '��{'Z�8�"���
pU�XdJm��4Hcw�&�v
����:�M����`P�O3���9|�-�Wϟ�?g��.�0��r�`i\*}����w_>K�����2��=����}Ҷ�����g3\ְ>�CYZ�^Jq���ɳiY9�S�Ғu��Yh������tj�Ȟ^ N1G��3^��JG���b.� ٴ�������b{ MG���C��+S�j� ���3X�~�k������5G!�*,�k'L��$B��R���v���u(��mG�`.�������a,�AUnGH��3l?#��u�M-�p���E��Yc�J�N<������o<��9�펗eO<},��^��W�Y���䣿���޴�ȡt�m����b�1W<pɌ�����7�*r"K�<�7Y��v�C���Z�w���Q�3�@X��n喅*th@�vz�S�Jx,���H�����~�}j�jD����YO�8�L K�������rc��/�k>�.c�K��vm��e$�:���K�E���1GEgf�X�3Y/#��QI���W~����`�wY�S`�삇ف������xH�/Bv��tg�c	eU,.�AE8�����m\Da2G�IǼ �Y�f�I��_�����HJl�쥾iR
X��9O���|��P�.Bأ������iS����"���]�WYF/�7��C�λ#{���2~|6�M�a�����lNWr/��M^�����h���-�k�e�e������iS�$z�|"���[���#NdI��Z�eŪ��K�ץ-�-���o�;��X{p�N G�A״?))k�F,�I1-�,9T��%K
�'4O��)6�P�p}�$�.�Ut����];5pF(�C�["G(����-��e���<�"e��<Ș�Cўbއel���h�'Ra� �J�fm2�ֱdx�.\��u_/�a��zIՐ�(��Cƈ|p77�r��ٗ��������n�)�~�m��L_��g��Ȓ>r@`_�.�����E��>�د%�����K��Fd��@"Ԍ����i���K�w�������o�š#�����?y6�4>�_�[�H��ҧ�Ջg�/�?R��	���gj.�A�ez�">&�RW+��>%d{�J�C`Ahy�4B�X锑)g_:"�n�l<!z��g�lS��-Eɾmh�*��	鐷A%�0x�ف�o�K�aC�C���o ��E��iym
ae���9) �u�8�M�6al��َl`��f<��#�u��X�?|gϞ���x�ĒA�T6��=`K���N��X�G~6;������2���7� �1�_59�}��U��H@�P^�Q���$c �2nn�(瀬���v��5<�)e{�q���A.�� Qjk�����f2�?�-_���t�b>�����[�Oɂ��{z�و�0_�H��;&�]�(��{l�r��St7��=�98���A��;\�1�M�r��f�z�zFv0'����9�a;J�^y_z��y� �U��]�DYa5;p�p:w�|:u�t���۲k�1������7�e�q8�Fh����w	�C"H�+9@���B1
x��C�o@��K�2W��mR�rdA��D�񑢦!M�v�*�̄c�^Qּ���M�>�h��?��@�Dz��n�,_�B���1�R�y�|dd$;~�x��=k\DK�NcH��!;��D�	�@YPpm5vqt�ga�Ɲ� 1�1$�
`���@DD����8�aE<��e��DB8Mz4�BF3E��UNX���ڴ�8�Ƌ�r�Ó��xL
��M5-�f�0	(�2�xc.�e�<䯼�gj��q��$��t��Ȫ�^�7�k��H2+��i���*QN�VW�܈ˆh��+�E=)�<�&��_�]�w���T{�_�@�12�ϛ�u��/�=z�.��r��%�U+�^+��^�*���2���^湥|�BK�(����kv��}�^Qo�k��o�{�g}x�\~+3��3��^e)���Em�?76�vu\����[�'4��h�c�j��c?h!����V��o]]w�9�E:1�X�q"-��Lץ�F�eG=�+ ]^.֭q�W��Ve w�;|���<�����3l��϶W����"Q�u�M�ҥi߁��s�MO��Y�� ���h�5�De���S���*�� u###�������|4�?t0���������-��~���;�@�I���@�A�o���F�p��8.��,�ۆ��B��fؠ�:����aۤ�_��O�����ңO�Ⱦy�T���/�s٧�����T�o�{�ڳNõ#Գ<;%d&�{������mi��-�@H���`9��`�Qq���[1�����|Z�n>�!��� !V`�і���ηB	ǌp��V�:l��Sz1RnL=XR�2�e��7/\I��~���Թ�;�����Dg�'�}�Pު�0�I�3n��c�B����	���"��	�[S�����z���ģ� �L�F𡱘~�6{����'�������t�ک���mi:��%
%��Ɇ�����\��I��
�桁� �/�F������ȟ)�R�cO��I:r�׻0�نi|f!��:�w{'�Y�jI6�0�2gh��	ed&���=-���H�w�d��kY�+ &��W@�PPku�%w&����u�:�0��;��O�����G����[_��b����x�n�e��Nd�w����ٿO��!�><���!�G%)�|ڽ��8�p`�9�@�	!�h�u�W���a�U��pq��4gΜq={�����*��D��Ȋ�<���:���� �}�ݵÑe���,e"kR����(o5���FFF��1�)�A��`�0'�Mć��\^@8�#Vst�*V=wb�><�fX�O�۶�S`��\�n��K�h|,��rvb�1tn���6`�A'F�o!���e,Q���9����T 6F�tE��l�gR��5��c���f��g��� �+(2%���)�O�Ee�R^E� 5i�\rixMx�`ʢ��L#����s��Q~�U|�{Ѧ������5Rqٰ�t�k9Dݣ�Q�(ߘ�ߊ���/��ȧ��F�O�2����ָ���7ն���V+��Wy{�<�^~�7�������~|A��x��*�(�����[1��2l`]:cֿ�?������b�R�c�y�z�`I����[;+j��>���j�@�D��P68�y�A�a�#���� ����(1O� �xG]9H�|aOI!�����@�bl��2E���Q�A��(Pc
&#��oĉ>)���I�iZ˧^ٕӧ�X��d}�ۡ� ײ�\'��� �Y5�Z`��^������~�Xz�� ��v(����~���ao���j�)��7! �$�(6���a�����E�-Ϯ}�te`�`�SO��p��������f�:�/����t��Q�0u�x�{�K��zuD����2'�8�m`#�v�z��w|w��;�2� �0�+��9e^`��zm�Sy�?EV��M��l���p��0h�̜q�n�!sf�:�̏��;N]=!σ�����r>�@�Wx�+�4�4\ܬoOZ���Z�D�j��b�t�b掭�xy�����&ad]ƶ#~�IBh<�2w���ߕ�=�8�F���������O������;^)�������v������O>R�t.�t�%�郔���o�~���KO=�D>|��lnR#����%Ȳ�D�T�Ƴs1Q�a;��}���2_h*����'�P��!�"�� �-ѭ��[�^ �RQ�A6�P�D�{h����Ï��\��qL��~��R>��8D�5�(���W��7T���R	��|�K_�O�>��Nz��A�@��iDM0���|��ǏòkE%̍n�*[�C泱�Ŵ��r�1ئs�_�2�o�ͱa�x�7�);u�s$���Ր��b�W����*A�}-�����Er24���x%(\�:��CVP���r����;O��ޠN=��c����x�C_���E��UP����1����x�
�
#�����@��m�HScғ�=#�!,p�p:�����
H?R�G;JL�&��)��6!�� ����dA`bL}P ��8O�f�b�"D���[<0@ @�\E������m8n�5����)��I�� ¢`��A �uN2����1�APx#�т,V �"�����H�E����0��M��;yr��֔/�S��փ1��5��'+�U�-�2m�5-�i�I|5k?yY�7�p�׽�Nw�@�^$��6�A�ۚ�a^e�����e����S6�_m����s�����V;$�G�0��h���V�G�MdYXLk3.ƔhQG[����uuΘo�(�T"��Q�����H峟�w�����W��L�����؅�)�V�綿 �RTDX��ڮ��\	�ڕaCH��E�Ɛ���	P[V�,ɠ`��ڂ� Ѐ���8l����k��-�����'7����|a��'7���s���<�u���LX���FN�<�cS#��!�98����2�����Bj��C��#5:8vbRy+�8�gG��sϫ�O~�~N�F�b���"���Lv��0#p½c�Y�`kf; �NlR�$���kDs%���lڍ����	������5�?���K�z�;�J:tx/r83�O�!X �P��WPooB�B�N��}��9=��`JINd�ӓ�>���|0�r�"�3l�,��3Rc"��R'*���g:-������R�ݤds�,�L$sV�d>�H��l����e�j�����)�A1�iCGd�{�����G�D�Vq<�����Gm C �&Ë�ڃ-���<責.6��a��k�NF�&Q �ԁ	ќ�w�N��_H?�O�I��?��4�Ӝ��{��?��4�E���|�������Op\0����_�����8Oϳdn�O���_M���(;wu*��w�j�E�>�,3A�pa4��T��5P��� ��`��@g܍����%l�u��3��i#jvf���n���|qj�9�GPs�h��`���(�OhT����{�A��zـ]v*�͗��m8��m��|CfG�l߾}�I�͏�J���Pj�Q�ZP1�_x��A=����r)7�䎃�������f+`r���۱�tۮ!�Akӳ+��kfjѺ���g�jQT섈�X�- �+��=X�YjR�����i�?P�������5�,^������qNU�)��D9k|[#�F�[�aٯt3G��Ѳ��#4=��Yɇ��&B�]��FR�י�� �kR��9b8.���nkvLȯAV�'8���:,F�P>x������ �LgN�# #	���� �CԚ����j	Hнa}	�~�Fr%0�%0
������R�$��>S��W��H3�\��B,����=����`�0BV��Dv�I@2u�l7�x���)��Os�4��/�1 P�\�,)
��T0�q�"#m��*2�vF%lA�z5�2#:a��r��p"L�Jpq�|��#]ď��J�ڧ�Њ(E�u��/z++W˨.����ž�Y}x���`gEz#n��h:}E��~�?��P�+�u�M�Z�j�������,�5����^�w�5M}�o�����n~^����b�;��4%���BA@�6ޑ��5B��1��1WݤY�6�@�\��;Eh<q:�̏���j�	��1����	1�/�2D��=�=6Q��2�S%�o�M���8�G�B��D��]���m���2In0n�]�=n.�Wr��֣��P��`c3�{����&�+�Η�,>|(��'R߶�l��>���z��ɞ;~��2�)w��z�̇�u���T�~ǠfR����ӓ?��桿	����9<����Wi�؋�;��=R��ȸ�`����i�i@���B�ɍ+ٯ}��3�i�M$9u�QP��*%! �B����s�CZ�
�]�i�>om� ׅ�oYf��D&u��ں�"�_��sv^�U�gg硴�|YڿO~�¥�3���#��Q8gl��F�A�
��=�L�G�/b�����l���i�e=����a~YV�+"a��K�(3�9�Ų�|���]o����o�����{v����sg��yU��=�������N?�L�'�q䗤�5���-W����˞z��4[�:ۇ��y�[y.�D�_�uh��5h������ը���/4��ى�Ysw_�B�mz��솃�Ĺg]WL��
x�NM�b��,{��	�mVwK�f���qm����95&�ş��_����f�6O�������\v�!۔��?�����Y�}��cG+�-�y�pv���Ʈb����ɌW���4ũK����}�����料��.��?��?s�b�Zt��>75;H�Z�cÁ�Z[ۯP1����Zla}�)w��6!`=�� r��zn�1���V�0)k]����q���S����i>}��n��uxJ�ܱ6�� 	RH���;I��mZ����|@}Z���O���dl(�D�.�]���A�]k�pTH@(����;�X�O�Om��"x�@�$�(����1�=Af����\c��<�JtY��ЌP7�`��o.0&`���t`�;�֥x&N��bC0"�,F�'
qA�<QG!C�R'�a���>�GU*�DS�%�Hr'�^T��Y�#P)�#�F��ƩW�cs΢��Gደ@�j�\��4�Z���[~)����
$�N1tJ��o�-ԥ+����	h!ѡN>��y��˯[�U���]f���f���"5�o�����K�/4B����bӣVF��}��lg�lB6�V�����>jD�k.�i���/kرj�}�;_��e�"M�q�����.��d����|}-���;!XO� Pq"@���\��@v*���@�U� ������q�D��W����A�`�/�EQ�.�o�����Ȇ��"@/N��kk�z�����!s��͘+����;m.��2��0˚P�w��݈��2cc༔�",pm�Tn*;@r<A['�b<�괈�<l�N��{���q	�o��c��tۭ7�ӧNfc����=��wE�jr�~��.�f��_��D=X���q>��8�sJͷ��&8��"or��������
gh�h6�w���ҏ��O�o��7�鶀��<O�]aB�
�����"͂T�YBwj�Z�DF����pM�6,�#��Q\�GvXD���|��a�!hD�kc���teā���iB�YH�^��'�0{�J���YoOf`����|#mX5���~�+Q/?�� ph��╳��]�Ab.'ķ�4u4�����Tj����^D�'���xnK;��Ɯ���`߬c�qfj"��[��Ỳ�}�S�#W���h�]�z=��cX_��>��v!0�?0��	���P�>��"����{өs�Y��:��S���*���,6��(�*��AP��G���<����2lL<,A�kˆ�����U����Φ(00U���<;���ƿ���w����3�Θ� !�����W�V˩{����2��t?b���;��u�^-\G~��7�m��k �_y�/|Tɋ�w�ȏ�h�#ص��
��Iys� ٿ;����`����g��������WF���8A�&]�N�p�3W�n�֫�Sn�玲�VϦ��gY�ʴ���W�6�t�M(\�1�^�|�2'���S(p�g}W�KEYw������(f���9�˱D'>��НMb�B�wˑ� D�6B� ?3Y�#^�]Q?{V�A���/a�����Ab&II@ɇ4�
U�n�v���x�v^D�Ote��Se]&�d�U���v!"s֋6YF� x�������9���l�ȋd�Wc�5u�x��8eu'�+�W핈W�Ǭ�/:����2��ȣ�c<�*�ތ�߫V~�7��.|�c}�����2jq�[��������v���'̺x��ʻau�#B�/�_p��×��˼��|��ɠL�5������T�w�� l�Wf��r���]�,s�q�:�\��U�YaH׷� �o|"3.).^�%R!˅�ZM��8�\A:<�F��H�iMy��q#���}Q�T�Yl�mQ��^Q��QNl�9`X�Nl6������	�gN���k�D�m�1y}���?�i쯌��7���&|Ϧ�^q'�1�s��qʾx){�}��ގ��e�ޖ�y�{8�R�H m����6��b�*���;�fsF��^XFnۖ�\D�	cI����B�goxӛ`���kBV�'�Z|�p�=�6A��XU��[�\�
�ϐٙ�������Fv����6)*T�v�o��D
�8�h!��D~�n��5F*�ky��6!�-E��2ZP����O g��!��}{_"�H4�1c�+��!L�����ƫ1� �����f 4K��+��\�`��r�8z)k�����f��]	y+Ȩr�p���]�xk���PZk��^�*��{��fo�W�p�r��w�˓Hv�:8�2�݂*K0:0Y1�g	��Ӛ�m��+p������3T�Y3���6)I�d[�BKVv��I�hbj.���K� �jz�S������A�1�n�._8�~�{H����t!e�����j�&`[?{�8l[��˲�E@��&�������ȁ�16��(�|wAX ]-����;�PTb_����9����׃�,�����a��{@� ���m�m�����]i�쩴��<?:�.@�Ҍ>�oKkk����:��׫�S�m�-����bi�<7R���.�F\ԫ�.�&��Ϸ�����k �$�=�zvb.��N��+�	��G9R�H�W�ߧ�pV�7Ď8iB����L@�Q����D?2�B@��+@�q��/P�i�Z�)��q(
�����(rF�!aH�Zd]KR{�C��A+�cS)6��@�h�.A�qEQ,[B�qR��^���.�-�  @ IDAT�H@�R�ԑ�V3��,�v����ț�5�rJ��8ի|��3�~���Kf�2~�ψ�e��4�&�ܫ�V���ȏ?�""�b/�/"��]��>�$n�V��ȯ.����F�W`�ŏ�z�K���终UA�!YD��Zy��h#���� *@տ����1�,���w��'D���S\E�����j�>V��2my/����o�=�)C$E���$+�o0���l��f��;��A�}��|���Y���� �Ʒ]">�R��k������\R����΋}��/�[�>'��*��-�G.	[�ĵO�K����� ם'y˷n��[WXא֑��TI��k�+ ]����|l��
�OW���L���9��Q��wxVď�֨}���*�kr>��;ڠL�xa%��֛o��|����a~mt	ĥ=�Ai@��	x�8 ��Fo�0����C�:HI{��T4�"��uAi��n��}���ȟ>�T��]�&�	>��5�����Ύ���c�f)"ɰ ��Z7�Tv��J ek3ykO��2�3���0e�����!��^۫��=�e
�k@
Dx�0��|��ڤ���-U��BV�#�#�u
I�J/B�8}�Ν:U�#}���?��P��/6��A���pAl�����rk6
�o������L�{�5��(f}G���>&�o���|a<{ͫ���n�rL�����z�Yi2�y�I�t�[�f���v����3 �){{�V^�t��cUMC����h?�B1��J�qǦy�t��v���A}���H�v�w,]�7�m�:�~�'mg�?����Lz��_C{�Gnޝ}�3��o��&����ܙ�3Xq��,@0�و�Q�o�	� ��F�*\�����-��9�c|�	����>�#�jiO=u<�!w�P��ꃚ�5�#�B������Eސ���f	��P���۳E���`��+ӳY6 ,�K��ŭ@�,��{s��2M}��z���Ş˼��|�{^/������0�������x��F�W��
�i��# d� ��T� <�o��(���D� j��&�B�y,�\~��$��K�O5����32��p�	Rp�� a#�B�)��E�J�7�����7OQ�2��FlD��퉸!�3 �	�g��j�2_^����5n��#�2y�w5r��>!�Q��)�AXī�U���"ylͻLSuk��]�q��TEx���Lc��Ri���=��~:�~�G�!��We,��2\|�8��H��u/�-�[�Y����o�y��2M�g�٢^L�j"����|�}� ��6���.;�|Dd$�N�#�T!RA�w*��R��y��J$5��Q���SaR����a|�6��H�`S�h'߽�n�/I� j _R���
��<�RY�uw��ODj�Ȑ��w*d���������.��mC;�@��l�!����3,�^F��16\Z�A��PL^�Gpb5[F>���h�00hZO�݆/�%��T�6���&N�x��0�ܖ�r�myj`�sϦ����@}Oh�\a���B�wNX�%��.� �G2��~m���t�:���/)`��h�Q�Q�[�ߐ:e�_eH��S+x�R	u�����؜9�
�OR����	̄V�Ӳd�tȴp��v��D=��o��巽,��׿����
��j�]ٝ�ݚ~��k�����{���l�������j�M�Jl�;���}?�����_~���UXb�h\�%�5�m�]ZW	jN�>��NgN�N���n���t��/������!��m1N�>�P���0� .M ׌���h����.X0C9��P�����OǞ~*۶}#�{�B���Ǳ�5�������P�Zҕk�Ӟ}�������q��8u�y���}��(���@.����O_�ʃp���d�z�M�T��\�2���r���U�-e=���0ʵ����S������O!������A��X��}�#�����X"���l�[*gXH���:Gt���v��HKX6Zt�r�����V�\�-��i{��e�w�i�pü�p���?����Oc���v�)O�91�R��=��e_}&�MMJ�F��1�XTO�溈ÏI�:�����$U�6@ѯ(/��gaȊ�i�\
4�Ņy��>�[�
`�3#b��ޫ�k7��l�C��a0)@	Ѱ[Q�\ѥ�b�p���n���������oPX�X]�a+�(�+��p�(M��fu�6=W���k�]d��<ˢ6�S�k�E�k�"�j�"g���*��dAP-�2{};6�-?X>����0cs���%�x,�M����cda7ƨ�wu�_��Q����U������+.A� S*�TJ#�Qq����@
�ζ�sD���w�A��=V�(�MW���Tm
q\���R�`F)6� X�F1��J�$v9�L 9�J����p� �P|�8��E����Z6R�?�Pe�5��,@��03.@	�//��	��G����5\�_�i�e�y���I�Y
p�3�K{��,��>OI���@�I�z�*�I�������r��͔!R��Aم���_��8��� ;�'�qO�_@�v���+�ˍZ#f �H�cfzk�=��CZ�U��Ҙ�l`+B���D�:}����x���W>�a������� ��2E�>T��4	p9�v6?4Q�F�Í�P�_Ə�Ա ��4*�3�ٿ�[G�a��e�u�Er�q�BE^�Auʗ���ٸ"���{͝�x�(),7r�m��Hy	$fG�w������{�Zv�¥�K��I��/�ϟ>��p$������K��ڱn܉9���/�#]��_�0\3�	�c7�'$om�̾�����A�1R���ET�GѬã-ү���WBV����H�ŧ�Uc[�`�Z؋�yG{%�>�T֍�F�ӥ������g&�њ;ø��7�v+Z_�iͿ(��<�o������Gqھ�M�驧�ͷ��>����󗯤_��_�d�>�dJ Qc�3�]7H���d_�ˏ����-��g��N�z����0����������ee�6�c�K�t�_�U��,�����R=�`�LD)Xm3�&��[ߚ�9N��E���}��-�A-[c�$�l.Q+
� �%�UE=�� �B�<�g�[��0��/Ӗ�����7��^���8�7���ӕ��y��e��ݸAI��=����&�5�iG@ ��w����s�
��(IC�lC��l�0VЁ�I"�q�� r�ʹr}�s}�N6��l�FX47ދx�_��E��4�Q6�`F5���=��p*�\l��<�?�^5<Z��dgT(�2X(�6��Ů($��h�_]�Q�(������"r�O� ������|mK�-�S�����G<��i|�N�x���?�v��T��|��[��w�����	���⏈R�t��Q7���2^�|���G}�ƠjptRĭFs�-��(�l"��{Y����-��e��7q���V�y/�և�Lը[�7��x�kHU��zu�{��Ҁ-+ +��H/QEV�/6������8�g�*l�3T��K�F���+ �}g%e���M�<�ؤ[T�*��1p"�f� ^K�����RzL(˿�$dC��놟_����MyKI�3������Ey;�>L��t���UU��a�N� T'^
�21�`��e?��&�b���Oѱ�
�N㳋�*��h�]8w
�؈��l.�h���A��^�n�q:l@]��^Ǹ���;�;y&��?~o�W?���쩧��%�Rj!�N�2j�m��q&I6�@^m��4�tx���d������H&��سc#�}�K�	���u؝�W\!�F�(T��#0>���� � ��|qV�O��<�O䋫������N�O�f� r�����3ڝ��_���Ӈ>d����'��û�N�����w��.(n���O<���F�Rz�d��
w3��[X�yF%+M���J���g�we��r�Hz�����>��5�A&=,:�����CٕKM�p�����"G+Pz�A��_�>l��������G��CnY3Hnkz��]�c?�Ϣ�S���'��v�ܛl߆&�<k�rh��h�uv�d�W��4sf V�$H��>�������}��ww���=s<��H����i��6�������i��+����9��kđ��s])�$�JU������w��]��Xj��f��ñ��M=�����C��e�
Q�s�TQX	�,8���f��������^,/�y��2o��X�2^}Z����!��j�E�/Y�>MG<ָ!}� ����6�V���"�5�o�k��ǂ��ΩHZTH�ѱH1�.��G��#�4o��?�������SQ��l&m�U�5���A��#������J��f~U� ����Z�����x~��Wd(~�i�Qc�H�|������$�f{#����lk��g���S��ڕa>Sd�>�:W?��g���^����gKy��l|3��Y_���U^_\�sĵ����&^��y־)���Z �q��'k?�<ծb�}-��H��t$�!Y�T�m��v�sHy� ��"��8�J��X˪�./��V�\F|A��P��q�{}x�U���hz�Q�K�*�埭,�b�b��4x7<�w ��k�E(L���
*ל�B���u=� ��M�z�y$7)�^h�t�oz�cT�V7])P��eS�8;��4��\�,7~m�HI��j1t�è��ʞ�p��d�%x��FͦΎ�H�������O��q���������cO�_��בqHSPo����ɫ�����3�ϤW���m{:�ܐ79s6;x�i�`?Fy�D (\E��r5�Ҏ�l�z-�,���Ԁ�ӣh9���хJ����)|ev�/~��K_�2,��lp���}6�0C����JAa�D�CA�����TP�ѱ-��S¥��A�* �+�^���Gf5]�Z�5D����E�,�lē�Ĭ)�;��D�����,�!F$���/W���g���n˞:�D:82c3���πD���w$� 6��6�c�\vM����顇J��?����A���P?Rz�ޕ>�_~/��faS��<�)��D1���[C�����#�M_��ײ����M�>��s�������miǁ,J��_I���JWN��w�o��%���׮O@!�љa{�x�Zz�g�Y�.<�=�P�?�?�{_}_�����t=N�������TzY��"����f�%��A���9����&\���|c����0q=*�]�����0]�\�_���bA�@|0� �L�i�M�Wv\��\*T���z��;��}<�p�\z���~�&��eCj���*P�u'��fS��Plm�b�G	� uz�E^����]���Y���o[��x��<�]��4[�4��c뷭�e�2����=�u�8}��$��\�ɑQ�SD�6X�~D#��kF�-E����!@<Y�p�Z$W���Rn�X�������q��_��x߰H�����k��B s���24o��<�@bӌ-P�
��.�c�U��؝�X�A5� ��-�m�$�"g7QИ���f��8E�ڷZ�D�?m
�����[ L���'b���lk}�Z�2������|����VMW�#^5��y�Tؖ���<����>�D�d����a���jċ��������V�,Y`s���o*�.n}�M�����^��&�"�]W��cN&Ex�q���aEw ���urj<�i � 	#���N�%�"�6>�2�k�t�w@�I���`���\醴|O�օ��&�v��� ��oj��݈�M!�1Y#������56
EH���v��X���7��#��,�%(K�(B��Î��c{��KO"g����u����~����ӕ�S	.�࡝�g�EchWz���ii
� -_y�ٴC~K�39���Q��V��,�ɍȹ�.6�S���pSkG���������`�]�Hs��ZZ��n,@z�a5��(�4c��~���E+�Wj�<dv ��l{�`h�L��|�q�'7I�_��YY��/��O#�-�����la�{��ӝg�B��+�0�|7�q�3X25���)����An����H���N���7�###���t�{�������z�;߉*<�5����}���X!_F��ܙ���n?K�.L��6�����b�+���i������uxj���U)=�ԉ����W�}/6��K���7��v�O|���6�_�m��Ϟ<� _tםG��v6k�c�6d��;�|�B�R��Qȳ��q����}�M��~���G������_G�#\̬w6��.�oE��j�c�9[�f�R ��W��`�3�����,ږ��A=��̗
j�۩/�f�O`�ADKD�u6�6��g��Ab!|�	cMȀ���b?d�s|���Ϝ9����G����{?�f��ۙo��s����ݒU� !�V�`�8�^� bo�]��sb��Z��O,f˰"F̡�7����^��z��W�����>���Ʃ��b�e��w�r D'cr �
�!�n˱e���x��ئ؍���Xdd��Bb3��sh̣�8z!� Ĵ�bD"!�Fo�8�c��h �.�݂�m\^tzt�Yb�*��?��s���a���sw��R1 ���e�H׀�]��b���ɗ2=Q�m�����"�ڙE#WYnq7����i���*�e� g�S)
#m����eY�7�ew�Ev>�C��|�UƲ�WV�7���m�Nƒ�R��^W~-�"�k�D��2"�?eXy7���[��O�Qħ�d�F����d\�\����"�6n���9�a̮h��pa��	k�<fH1�����/(X$���\�[�?r~���cm�TR`�?��s���yI����]��ĄJD�؀=<V� !�����֪��|�v;c!��և�^5�ϊ�~�H�j�X {���G�e�ٟ"\"3R�dm���m�X��λe���0���2K����"^#l�[L[2��@�']�Z�����ƛ�!N����l�~������ܱ���5��A$ֲ������I�h��ut�g篎��T��kj:���.�#/�\D����`ؘ�t(ż�@�_��܈\���؞���ԅ�5�Ti䦧o;�LV+}��R��ϟ���u�"ٸ[�����G�v*���������+�Ԃ�;�Mt��,�h���0��ؠ���H�֜u���}��|�+i���_=-3_Xi����3��c�1�F����a���;ƺy��]u��$[t:���!(�����O�="L�g�_��_O��!@?EN
��3�Ҟ������ϲ�������n��t~tI�3\�Hc��Q���aq����я�nz�?yojކ���c�{~�8��̾��G�-7߀UH���J�z���
�g>,dhz#D�������4r����3'�G4��w_����aҌb1�7úUz�_K���*D�3g΅�C�f��oqWӉ�3B�sB�#7ߘ=s웡Xp�̙u��W���ޖ�?q"��h1���$�L.�+��<d0�@d�IB-tw��逢%���m�?���RVg�;\��(���
������T%a�sDJ�b�'�1�X��cS@6�Y#3	���E�ΏM�a\�6�m}ߔ��R�/�\������2��򶾗���˼��oKA�g�hn�7�O'��Ә��!Z������vp�FFFҫn�%kC>`ABA��p�jq�K�YV�yq�<3s@�b8���M�T� 	+�����1)�0L#N>~�m������r�(A�����#�����ƎL��(����*�5�ŘEdI6巨}z�GRXE�uy�d�ү(�,�z/`Z5��[�җ�J��օ�n�Z�`�L/Y~5iYFy7�|�{�i5����Qˊ���q�ߪ�-�^P>�,8u�IU����fZQd�ү��>�9h������|}A�����~Ɠ]fINL�������#��}mqc�E.��(�Z�<���1�)�"B#��l��[�5}K!X��*"���b�G�
J}W;p�Dᦠ:�UY�ꊱ��/ɲ�S����DǍ��i�����q����Fk���l2'!�����L��?���l�Jv�c�zZY�wu�/~y��L�ڋF�ݻ�� ���𸺰�Ӌ�G�>��P0������]�pH�w�����l��w�X�κ��=nJ�E�0���4��@Z���sօ4�ɧ�;�5�߳rZ�P�i9iinB���l=��!^
�+�Ĩ�0��"2[�<7��(��G�;�l�;�b��1ޫP?�O�`�0��@�#<c��p����G��7�%�p�p�ƻx��j��н;�T�����`;�|V�*Cx����D���\i��#tܞ��1�Wa{v��|���_?~"�3&�DքY�&�D�;�VpS"ۢ!�_������06�nD�PP�cp8(mX,׾u��%E�q���PngyÜ�]{{"��.e�_��D�u��K��v�6������@�����b<r֏,G�S�x<����|;T��CF�٧�f###,�)˷�(��y��'�@�k n��$$�[� ��ڜ��꾮�U��k׮�����Â�J����9)08HN(��3104�Z_��U]p�|=H��cD��t�c[{3&ث���Y�W���S��g��7��^e�2�|/���WƩ���_,�ּ�ӕ�?�3BbC6 �o�*H�<���r^Y��>&R����
��=�w{�)�`������������I�'����H`����ΰ?�X�sV�/NN��(&w����:h�a�j��9�U�^���ص ���8~e&��O|1��S�um[x6�G�ĵ|�>a-�i�������8i�a�8O�k��$)\ 4T�y��Z*���ʔ��T�X �h��;��3���Qn�����F �R����(Eԋ�ZE��;���E�~��5�p�Q�P��%*_���$�����Op��1��!�B�#�y �S���[���szF�K�b��K���Q�d�#K�/�R ��l�Տ(��(K��bĮ���ԻO���Bk���i�n�"��+�9ؽ�h�@����hE{�L�X|a]ؓ<�����0XF1����� `��N��Ņ��D�j�������붫�sIG���BEy�B����KW����)	=�{U{��j?�VU}68��~맺���p4��q��\�8�42���E�p�Єww5{D�[\�ͅ�-e�l-ס�FVRb�8פ��/��g�� �Κ��L���Lc�� �1O<�ٚ���L̈��k�+���	Z�n��5��:�+83�p&���#YX��\�k�(����{�S����E��>��s�f�ǝ��I�tjy���_֯!���8�e�d�fc�I�/#|=���|���LÃ��Op��MVf�u$��E����D�*P�+�߮>:`C[�t�,kwn}1�@��(J>;� ����Y+2_�+��s'���k������7w�|Z�:߃��4	�~a�A\J�cKl����s��u��+�뇇;*�X��@xް4���z��H�3�]A�H�r�fj� <�F��عA����9���l����D���Z.K�bl�Y,T��&%P���+�����43�Xd���П�`~���pD�s�^����� �6ء�0�ֱ��۞�t|�k�ͻ:���ѱ�~�?����J��[n��؝z�b0��2�1��{c���ݎ�˸s[�uKcv�����ld�m��5�_]������2���\Ϯ]9�v�ɞ���k�_����|7�ɶl��]����Q4����~��6LD̯���q�]�,�·�� i�H��v����o[��ߵ-�Y��V�!BLг+���B����ߝ�!�591�N�:�>����pŚY
�y�,47�+:��?|���y��D>�q�d��C�]�#�ʃ_勧�|*;�����o���ۑ�����T��K+�lM��?���.Ⱥ�s��o��S����ԕ��3����!�Q�8�D���>܉�U~���p�^��/�y//���a����l���[Y���F)5,J�:Ŧh�{[4��	ع�â�� Lέf}� q{!�M��x�j�0���\��v[h�*͑~3���i;��C�w7p�;Rܳ
^���Z�}硔=���t�᧳�~rn�n)^�M{��b�ΈA���#��?��k��T�e#n�-��=jk+��î!��F�FXl=�E�j"�DՋ�"��)�m��i<W|SSF䈢��P�jQ��=m�B����X���{��">��V�j�ti<����2�RS��|O��t��<,����i�I����&��"��aY�B����T,��� =�qZT3Vm��!�H!�����@&O���j�Q�VfB�7j�/�Yws�$�y+R�R�_�m���.�e���/Cbz��m#t�S}>�g��6+�=L�}�&�C�S�A���@�";�t�d�x���D ,�$�e�r�����.��Ώ�x毌�T"�u�a�,�8\Q�R!FC�":Z��.��=��֟�t-�g���P�	�-P���6��9n�����T�n�=�OL��Ξ;�@�dȖ�66r5�._��|�Ԍ�c>� �5(<���)���C�^H;�f��q�z9���hl��u-)뇅㬫�y4�~:p�2��q��.5����m�P��luYZ �Z\�N��ar.�o|�+#ߐ�����P��=8��ȕ!�&��x@�P&��T�l�z�U�C�����F_�.x�[̱��Zq�؜�/�9��͹�Y[��ǵq��&E)�@�<�Hv��gӮ�NWQ�0lay����l�����̉�y[{g�[�ĉ����.ܰ@1`�3]�t15t��N�>�z�ѿ�Z����@� P �N9�3��eCP/_��]���\<�����i�db�$�$����:��_�!)5@Y�'��g��uҜR{¡���K�;�� U'�7`����{�o�g��p��,�6p��?�lA �k98��d�*~K7�}��"7h&B��R:��C*l5�#�J��>T�72��C�L���C�kP���)PR�p�2kjxxй���o�V��˯=8i����6���Wl�� /W��`E�ȸ�Ա�S8緝�܊��^[ߍ[�o�	��V�-X�����k��ߖW}�2nyo�������������<t`Lf4��J���k�r�*[�䴭�΢[������$1$�V�$D��;�^�at���/�A�e��;��e@k2��j��.��K���[�ͺ�u�a޻8]�1I9Q3���̫��8�G���*�P��[�=�T1��hC��(<��D��5��!ň2��R9��8n@�IᮥڗEH�(��=ʷ0������o����I������{
Z��ĀL7��F�La�muj<���.�%5A�zzӸ� ��0ʫ��!/Y~�T�O��^14�OpsAK 6o<*#�Q��>[�˅�ԓ����Ɯ�)/1ۊ�Rv JAq2�+=U�n�����BP�3:�kS�j+��Ѡz�8�&�LX\��:xD	 X����6v�;s��Z��X�e�U}��(�-��g��0ߋ��TT��V6�G|�eύ܉���Y�c��@�E6�i���i� �i�TM�D\�0m5�
�΅�k���b9����2#�@��]�(�oeHeHu0�C�<�YE��X;������egg7>t�*g��&��`�Y.�S �8s��H�z篲U�=�Y?�ݶ!Б�|���[l	��]lb=}�j��i� ��. �8p(ol�bJ3_}��9*S�ښ���� n��Fp6S��M��;z۳�I�-t�5A])Ɣ.M(�E��9�A��ցQl6X|�M��鞁���&^�~�~ｯ��]��N<y5���{䉴26�5c��҅��:2&/{ŝ�'r������|�5*R(��T=�%�U�.XnjS��1���LtOo^��y�Ǆ N�W���cC�~�?~�I�e'������h����<���oH��M���Nb"a5��Ȱ��q���<��w��{��w ��/��+���/����_z��l��[��'��kNg�=�z�Zi#ma~aE:=�������&?t�H��7LW&.b��)��0�����-I�1Q><�G�@p7S�V�wf8�mX��n�H-�1S�h��oo�,�8sh[z��c����6�V�<ujw-��'����h�/��Mx��^AP|(�`�`�+ǎC١W$�U�Ư����i�'����D��D�����ɥ��b[�rm��7Y_qķY�ϩ鱀�M�T���Ju
��dn��K�@! �-Xذ�y��k5�c���|ny�y�tI{�?�D\���K���� �����[�e�ͣ�\�W^�����[gs`��V�0��UA�040P�@�������'_Lo������*�����Oj��A�d[D=YЇ.N��1l' +<15�EN�&�!JUCFm��"�z��8�U#��S����]*]�& >|^�D�.onD���B]��P��HI���o�e}�+��lL�p�e�|�4�rE���Z9<}:�Q�R��#J��#a��J1#Ҙa�2a�ܺ{�Ũ0$�Ӗ��"Kz�>]Z>��D�#�Mm��u67Ƌ�>�i�ȲNEFQgr٩^e�!�>� �$HV=-(���_4�h��p��l�T�]tQ�o��l?{��jWkS aN�n�/[������K�Z���8̀Mh�ڍ��(j�ΜКK�Z}h?��D���U���8E0�O��m���c�U�ևT�[��q���m�+�bM�&AlaN���f�-�2���T2Y]\�k��s9���M��ȉ� ;��,Ն��jc��ǲ�J5�X=l`���"~��a��oo u�S�'a(wAeP���g�Sʔw�F����M�����vݦ�Q�����´�^ݢ�M��L�#�bM�A��[��[	���CuR�|�gD���a�e��cm:�U�07��Og��B:�[�^dd�a=��r����*����~���G�8����'��ӗ.g;�w���m��1� U�չ���i�Ρ�����(�};ve��_�x�������V�1/Б�^�������,*8�l�u�($�F�V�ؐ]&�誗���4�S/�)t*�Qg��/���c6|x��|hxOv�����W`��:\�6��}=��v<����?���t_���<�>�[����q`�>��1�|;u�|���?����7�h�~�vZ��P���ξ� C�VRwGz��SI���ߗ_� �<m��փɆΞ��'a���R�T|Y��3�412p$�`���.-�V��P�v�����ęG�y�|����/�xdO=��Д<s�2?���#W��A���oۖ�p�Hv��s�����������N���-(bՙ��a�"��#����ȳ���YR~�m��|�����ӥ�W��K�sױ��a �"a���^�?y{�ˮ��w����X�J*Ie"�$b E������~�>y���-�(2�29 *��4$!�SI����������9�nU���ޮ��9g���k����k�əg�W���U�+Ի[־�,h'
�j\�Gΰ���ffb'��%d#�$U8�!�xtP6��ޫ8�@g&���U�W�ճ!�Ăi�M�7#����j�:���;�B� ��񱴀�|/�{;V{�O��;�W�~W��m��M3�>De#�z�S���էD��&�{<h���)A�@�b8EŎ����9���BH	�:��*�+���ү����ŷ\�,U�8��ƑG�jk���Y�>�@-����9yL�/$��ǂ���^�l�J)�1��J�b��w��C�S�1"eE|�D���U.O���O`�Q�_��;'�@g���W�-�S� !n�F�	��9��&v�7`������a�/��Y��Q����	��P~hL�v(n��N�������:Q-(�c�)��Z�Eǐ���pe�����p:�(���f����[k��\f[����m$���@��%�X���O��(gcs毞�q��yʩX�"�F[��փ�uS=�� �sUG�󉷂_F�W�������#�Dpk:;{��;6q&M�O�ݙ���붥A8�}��*���Lk,"��ʘ{����s�c�Z�"9�_ \�Vj�_�s��.�KIT��[+;M?��iA�(f��76c�DZƋ������t��/�G>.�n����n��SN�SgΦp��?�?������r��K/����N��2��XgK����wC��?�X��<�`Q�$֓����Fr.�z���D5\Hzj*��M�#q������s���v����q���aS�vҗ���O��g�u'J_�S��4��Sp�WG�'kS����eYO`��������N����_�;p0_G��{%Ðe�a�`۹<�����?K��n��,g]��E"N���_�c	��)%�D��w�[�?0��_Br��b��H� �?�G
�*?�O�����C�7�����6=���g��5[��c�O�vu����=����߸����cr#�i�k�>�>��}��.�]H#�6�6Ph�r�4yf6}��_��}��40ܕ]�s�9�����97���KnLm�������o�$�
u�e�XbC�0+��Χ��i˦n8>Q6�,��!���ġ׶_|i��?��W����v��1�i�����q����f&��J�i{��{PUj���u��[��ĥ��<��e1��4p�N���L�-�ܒ��ߟ;q4�f�Xlt�1��|�3�Ⰳ��M�q|N����7�1bkŸƤu��Xρs�R�s�Oz��N��m/�Y�b{4�_����@���^��Q����_�������W~���Z~3[AL�uB����r�Q@�u2H��U ���i����x��\����t�E��C�iI]r�SO\�+�mA���ds�:y���a�ƘԿ�#��>��:��M�S��2�wW��yt�Q�Ȥ�:iۘ$���\5��6���Pn��Q�o�˺����=�³����_���|��v����?z	�>���O���t���UO��/.�JP>�L�^�v����@�R�޲\i�W>t�3޾#D\P��9���T����z��*���zZ�z�b��J&��1�ۄI�ڭ��p�r��i�I���m21�����l�߀ �%C�s��!!g�pW���mv� �B���\�qiJjb��NG��SpԶ^<�6��h��j����e}ë�1���;~G�����jHR�ߍ�v[�zp8c��O�y"�m�/u��~m)����jOB��㧎y�1�o�d�I	�������_�-��	�n��"E��3�V�yD��qapL���|Fy>%r���7� ?.%�h$����NSׅ�^�:M� �9�~N����e���ze�;mF���]�{9AEV�w]��Qܹsg�ַ��P�Һ���).G�Ћl�Ť�#�؟~*��]���~�����7���۲�޾|�G����^�ڈ�fƱ��gi�?�|�D�9p1�i�\��ԁh��k6�����X��u$9;���SY?�/�X�F��8��Φ��̴����=�fH��o}Az��r��l*{�sn�ZuO�/~��|Q��ZD/�J�m�զ�N��~�s�o���h��������cʆ/,��ߘa�8��7�\�g�W��6��A������x���=��fNZ��b�Sl���rY����n�S4��V�>����4��q���-%*��ږ��������i��u�\yґ=���a��M>v�y�lW���r�"K<0M,3�ьy�;��:��{�id������|~���nOo���t��#(k�L�[�!��C8?��f�϶&4�]+H��  @ IDAT�:!x��I�cq���t�� 5�x��Q����	�r{�/EA����8������oE�1w�)8�����qR���a�:-����)s'6p�`G ����@zZ9��+�S�C�pReN0<��@Z�k=|�6.|V�a�7��]�*����w�[�Uq/|V������w��~��y����/����Q�� @�m܆�?'��;>5��	�yK��	�IQdִ(�,z����}��j���vY�b��,�1t��%-3$v;�����r̵|���s]�<5�e� ����l�#�I�Y�0Š�b!u.c�(K�����V����Y�[@DB	����fHI��RF<�>�뾴��ƾT��/���FҢ?�^/���:V��_���KO�Ho�a��u@��hQV�;T��4M/AyzrH�pc?W9�ϡtȮ��0�˯��bq� ����P~������X�y���A.ѹ��Qn���m��70�bI�%v7Q>��ǴO*�H�hA�B�8`�].蠥��B2���]��u�jǸ����G%�k ���E�9�bq _[d������c�DUeX�!�Sȋ� *QLX�M|�w�1�xU�"B�9�"���άh''�����pO�k��9B�7��;M�� �l�D��uY"9�I�����~KdR�u�Jp�/!C��+jaa �9�_�����2��*X��fl�\ː���"Dt*�����(�.�>�!��S, ��S�G1Hk��1��,7lق.�l#����
� E�:f��;5��8g��W��e��6�=�����7�w��=�&��4��oI?�ӯJ7>����/=7{����~��?)}�ٻ��>v���b��W�4�������Yv�3��>���f����{� �N�+3X�;�q.%]�K2�i���' d���/���f߼��yW�lv���\�r$��-�	�j1��?}>�}٥���S�/\��,Z��!c�Y�(��vLJ�*�*�����þ��qU<���c��(�R
��^�}��]NsWWOpה3`�)��4�ɑ��5W_�ӗ=}
@ZɖXgZZf�$1vXD������?�b��� ?1���[N0U����)La��F3�ί߰���d5?rj2�sOܖ�[�?��ǳ�S�Ik���NP���_3��d�Q\}tӢm�WP���Q��¡ۙcN&;�����Y����Աܓc�:��l���c4� kl�dDw!6c��b�6�U�]����a�t�s���h?"]�[Z�Op�Ob& �Hr@ �8
C�&�6��fh��K��:����}�_^ �k+��:�f40O�~6ud���Ɛ/!2�l-�Gg{6�ۭ�NH)E(��V�O���K��Qa�'Ʈ�\R�q����)�1�����|D���#m$eX�v_W���qM؛�ޫН�fs�[3|'Q7N/�4/�d�.���J���@������@�&㐑�X#=YP�%����o�]\i�f4��AҖ̀���� �ʶr����T��,&���z֫ʼz�<�ix��T��*I�H~X����}�Y	�FuP�!3&� c��zc[���w]c���Eh���Կmo�����ӿ��X-@L�w�]��v@F�:x�d;��8���J�wE.Qj��y�E@C�K,���lk�Dy�  ;H'7pGJ��%�A�a͖��)�*_����w�������D2�dJGO7�%�)'I���:���W�&DE\��N��:�g��OV��/���}a����\eR}Wy�lLax��,�-��'�!��ɢ|�����v���-�C�%w����]mE��'m�3�eoEm�;6���i�X�2�I$I ��N�������1��p�ǸQ>����2N��g΋yV���o��ᆷ�4���C|m\��Ex���5K �Ҝ�C���ڝ�+�ba�x���ԅ%�Çbi|B=���-q�=�x�E���������fw������g�{r�SM�KgZ��zNv�=����#}䯿�1������;�[Z��<�`����+^�N�Q_����|�;Ր�U�z���C��nDv�����UtI��鉴2=��Ad?�����/�4�{�W�=�_C�}�C�ֶ������d�a��[��βɕk`�1V����c<j5O2��/^/��_-p�F��;v�T��$�#G0� ��������d���aYzKΩ���������96\=�=�<�BD}������o�@��+^�Du���1u��j��M��� ���y���f:�#�ؒB?i"�-_^l��֧���\���g����V��)�|f]��;A08�
!;������nLC�3�w�r�I1������ܟ�m� ,b׊y$'�z�5��b��B����p�~#�#!د�t[v�����-,`�u�)jC?���J >�:��9b.�=��@���L��9ߜ�̙�o~�7��|��+0T�4N%:�Т�F�s�'�ĺ�:����/��2�LA���p��`����&��w�Wũ'�ż�Y@�����G�͘b�v�]��i��$�m��Q�2� D�t:lH	�`)Bͫ ('�-K-Vt6�r����b!-[;IiM��)Y��C�DсrrH<ıs'���E���"�E�M���ͮ�x�+�.�s	V<�}�K^��D2�v��v�9GN7� p�W��uϑ�"*�GIlDذM�����'��"n�fA� ��B�Ά�Y@����qe��@Q�Y�n�l���h0�;p\���U��z�^��N��ދ�z�l�;=헅�玢bamx�ػn��E
���lv�P��4�Tf}�vLU^�^}G��4zB���S�������3����c���眲(�)���Ogt�k�
r�9�(.�Ʊ{=�)�8d4�A�S(k<u=�23��@#��s۽���XX��Y����Ɗy-����mؓEG��'�q���_�#�S4��N�>���@�6�z��E��	�>ʇ��a�st2 ��kǝ��	_a>��>1˕�����a#�i�|��a®~��BqT�
���y2̣�������*ӛ9�#O�o%q�N8�
3�A�XV0a�pN��^�81���;@z,�K�1�[�mC�'�ߐ�lۊnљ��Y��ޙW��r
SJ���+��ۆ�p�*e;�N���҇>����?5�t�[��@ U��t1כ�H�'�����<�~��0F7o˶\~i6�ܖ�Н���,��U��^�ʓ���}���<����A����_�ŴeXN�����0�5��ί�6������������lL?���c��������]�>�����WD0�4gXtl��fqg��E����iy�����)׈��B���\�uf`@�q	���o7��*�۸~0��=�c�1{�k~<۰q�G�i�q@���X&Q��`,�8h�OE{Ζ#�8C�{C�H��td��\�f�M2�LrS/��ٓ|�$�m�^���3�n����l|���D����مM����Ԇ"����T�[�E���S� ����#�C�轏�h�c?�:����Z��#�F僞�=��}y��Z�09�m�IlO�h��	��
	@���h�qQ[��p�������[B�{��n�p9?mGj�1)����_\|���=�X<1A?IȺ��,Kt�x��2Bv�H/�3ȡ٣���*�1�61>� `���:F�����+���g��~b>�f�2� :=J�d�0�Ux�w���\��Mm��C6�|Ttm�����Ho��2�~� '���u����oY�w�HdOT�!1������0�u�_��w��e�P�LP�"*��M�f��ՒɈp��v e����A$�㩘�Q�<؄�5����Bg�)5 �����@�L���ґ�E���/<b �/^"�._��=!�9�o�2M�YN��||����
5~^��,Q~Ywêv��Ţ[�+�*@2�u�@|t�
8��J�ru��q.b���y�7�\X_���?ZS�����X� �xT�����.��&�ԧ*��^×`ǻ���wSH@�K�ّw7��S�<� �c��WDx%��D ` ~C������Xf�{����֘�iK�JW=Mc�x��Db��Y��(���%�6��A� ��/�c�i�]vY�m�/��$x�#8�J��H|��\h$�pQ���8�W����q�wRh|����W~�+�7��t.Q����S��X�ҢԳ��i^n�=��ndUw��p<v/ǹg�4y��c��/�MTg	����3؉)Dz�gg�;��V�R(V�!znV�C+xm	���}g��zy�ko��X�^ל}����1�����4�z*?��@pO�1�ގ��GKmH�dǖ�k_y ��ze��W� ����^z��`���!l��E�u���w���L�_~yz��_�~��t�}������h����`l��k����D-1����ؿ�{���S���X	g�B���'�s�k5ۺic�%8$�ҍ�ؖ=���&8�!BO\Ŗ������R�K����'!Z�!N�ft���D����;f'���;�e�4����k�N�ןx�O��镼�m���;;v��������3ci��Mi.���N�����D+w�9ぅ8���>������+g+�qO Dv��|�կL�1 �<;�x��p0�053��ܵ%��e/�9@�	�cG�y���w�6��pEYݜr�ƙ�����ԉNbø�v߾}�g�������mݽ]!f�kj�;�νk��F�)�򗿌N$0cn��M
���؜�Ҟ��dwwg6�ȮX�(8R��1 �DWl5���0F\���!�i��b�����>(K f,���������=Yz��9טg��.,�1�0(����Ѥ�̂�"7O�`����ʅ]@H�VAB�)V`�Րg��(J�^�[���@{���Fq���Ť�Ol��'���j�+΃�Cv@�Pى6C���$w���c\��W8�&7k��bj�,XL���f�F�+�JV�"B�F�HS��]�+��s`������G�}��>�/��2����?�CvV��Ox�U=���ʯz^P|=kj>ƫ����MŒJ�>����d8}^��cX��z����_UN���T�;QCB,�8�ZҘ��-�?V]��.] ��|*�h(�� �Fk�7J����c�Pb;Pl�0@�x�9��:7�B :�<@�u'��0	((�*?{�w�T~ƭ�U�t�Z��"B�/	��U�V��G�Kh)E	�	Oa������|���ʁ>E�\D�*:�r�h� ��qg���p1-�����rl���q��tc�n7ƇȦ������Ҫ��q�wy+�)h*�	GҲ���,�i�e=}Y�8��VKk�8ݵ�Fgڻ�H-��r!%���j�I;_�ƨ�\~r�u�3"E���>(m���&1�����	�ڠ�I?3����d+�H��0,s�5�6-f�����ߜ�卯�siMs�������R�����Ϣ�Ҍ}��M��@x�H��6(���9����[�՗�J���"���>�I9}9��]�=?��_~,;������|��qw��eig�Ά׮�3ҍX�4�j�J�/qH'GZ��~6�8:&�/Ɖ�C#�*X+����_�K���,��c���M�sL��'�K^x+���Z�В��=��F,�F	�2lYu����i��
mpt��O'.���D`)k�#��@k~dz4C�+��,�.����78ѐ1�B��E���6��8��F`Q�j��~y��MD�T� �
R�7gd2fO��&(�{�d�wnO�B�� �S)۱c��d��%����0<�/�Mg��б� �� "HI_��!���b�	�uΓ����E��M'��9�z��Ӵ�vO9]pX��Eq<�I�xI�M��s�bO�y>59ż�Pd�!��fA��c���nC�as��md
�.�������
�a��k|o�[�WO�b�6Q����*r<�oc��{c���*���*�*쁲�T!�x*��2�#��CHS��Eյ�j��r$�O+
� |���?t6�ƙ�PA�qDHL�B�nkbM�z菂�!� #,�+.�<h�f04�� v �V�_�I<���6]p����u���kmaj�a".�����O�:Q�9܍�3�H\fQd�_1�'�0�2�z��u���>�q� =�X�_�^�o��Jb�P����9�-?�� �|	��L���U�]���'���«g�ܷ��P0@�d�"����q\�$�P?~~��YveٮȟwG�2��g���2��Z�`5�Y����fZ3���P�#bR�(���aeIц(�軲����cD����{�����ֽ�����s�6�|��M4L�n_�TdE��=U���mCd"8w��enk�ƅ"�Cp�$<�[�"�ȃqT�&�����_�>����0�H�/"��2�_|�4�M�v��чQ�8?�"��2��3�pd:v�8�gE����At���kԳ˹�N��B��R��!W�u�B�AbAV��������iǶ]<
i������U/I�;o�Ōu>��ү�/}��H�.�6�ͮf�
'7"�ڼ5?z� ��ڸsl�Ng3u�^��7����_�=}�wA���k��p*f�W��tC�˿�_������o.�:,�w\�/r�p�S}��#a�6�U�K��9\� �a����Aa�/Q �J�D8��|jz)ۿo_60����+�����?I��݇��l�e��b}��!Dty��1�ͣ�������m�J7=�Y٩�gӽ>�ǭ
]���VTp}�������x�E"p�c��p!���� �.$t1N����m]pWh�I�qʿX�Y^��eǎ��}}�
�b���P	 P��[#����.��9����L7Q��v��dc�Kن�-�o���	��6l�Da����4�4D��I�H\%�>�V��sv�ĒP�H���.���c�Q�e�p�W�,��O��Ϝ�/�� ��o�!�#�����^}�Y��6D�\�ÝE0��6�Y�J��g�8��}qj:[�K�aGn��|M�h��>��rG���Yw~W0taX=R��n��o�D�����OU�q�*�_S��A�?��O�4� P�PkC7��(� �3g)��!h��A���j3��@<�f��3b�
2�b7[=1j�s߲�8�?�-�A.�Q��fS��)��࠿�Ht��`Re{��N����wdg�s��3���h:Ii��4{�-�\����<ə^dQtLh:���"NB������ @{�O�f_ֲ؈Cx�"���g�_���|�g��Ti��#&$���9�d���+������'�o�|-Ӑ_�8�ǖ)��*�]��>+�>)�t^����0��gI�TM����������\>KV�k���<��0;�	Ģ�-�7�S�H����;�& 
���|���".���40|�8!3������-AÙOYN�?�ddF�F��U�x��)��13� 4�9�S�%�X���W��5Z�CuJ���\ɀ�"�����UR*���W��(�A!D �ޠD�f�Fz�(\�E�Q"v�*�(�9KD.��s7�բ�� ʋ�u��W�j�#�}c�M���ERE�v�v]Hy�����߸��vvϓ�?215�FOτ��S_�DÖ��d6��?z޺���I��?LA88P�X`{~|d<��sU>����n�p���u���Si�Tk���(J�/{񋳷��O%� �j·��G����3i�u7a:Qʷ�g��m�}��@��47~��M��Kwl�.ڴ6��`������;m��׳�N���
N�=p�7�Sǎ����('9�����c�y�t��ٸ��1/�k��Ⴉg����_�?=����N\��/�9'\e��` ���-֥������?s��6g���7��M���|z��Aڶcg��ݮ�2�8y�3O �ð����&6��ٮ��0?�>�я��}
�⋾7����]��O~Z;_ywWq��d>����#����Ox@Y=�b��1�w+���$�0_\qSkͻz�������2D�ԙ��#�V�c']c�6�^���Sܯ��X����ɉ���Z<�i<�<�� �ӑg��r;'䶫��n�t�D��)q��r bcõ��z�-� Uu���½���0��v��.�o~����tW4v����O#~��c�AeZ	#��xL"���g_���_��ߧ���l���4v�L��5�8p!�#9j�Ev�	�ݽeS֓�����c�����۶���1�\��z"�$�<�#���ر�o��?������8>���4�몰������?*�-�؁�A'G���]����Y@:?�67�p�ϾiVK��.QDخ�L�V�#��P� c�5!���25�I"9w:��
�����`Ec�� S,Zf7/�g`�b�3nE��}�Y�٩+��A�xR���u�A��� �ͶN�^۬G�t�r�#��L��_���B���#jC�ʿ��;�F�e���'K�W�$B��QU��7.�/���,lh��Ic�IY�
�Z�Q�B����/��#%���yF�~0V]h��9� �Hm�*��.��\���Z=��8!��C�q�fY�it|���q�0"~A �-@���O��+�(�l��ˮ�wi";�/��U�����#ލG��p�WI�d�ښQl��݇����ıc�P�]Y�����{�惜߭����Z�}����;��S�C(�"!%p����ȸ8�	#Jĉ�}��-GW�i\�Lk�]�3Һ];G�X�0�"*�k(�B��.��˦NX�ю��Y6z�,��QF��4'�:;Z�t�C���)G����i�׆����4rx/vT�����4������e�vw�����I߼�!��,]�kgz��~
�F>�t��w���?�������}xsvx�l]�p�+�U>3v����S��^Dvߺ���~��4���߾��������n�_��y��0|��7�>f?��呑��*��c��B�K�Wj��j���!��"���g��1��ó�ST�[agEf���?�9�A�vuw���H�����W~�W������^����C�����'�0;3�^󃯅�с����?����?y��ʿ�y7��\r��i������U��]�l���8����y�o�`%����Վ�Ls}ˡ�����G1�0�}��?�Ϣ��gj��-V�Չ{>�B�������&}��X�kX����^�L�,M�ѳ��ݱA�agK����������Z����8�1°iv�;�i�<ͱ�m�|�ۍ���횺W��88�{j�ϼ���g?�MG�Z%�<	'�i��푏zK��*\Sw����S�f\�c�w��ɺ�����dϹ��������y�ˮts��k�d;�|#�+7pQ^wsvtn?�t��Y�0�\�Zc��3�.�=�*��m��m��5��"��`�q!N�PJ_я���ۊT@4F�|��[ ��U�|y��I*�
�K56�S��_�HiWq�
F6l�t�mj p��kU����z�:J_�5�3��R]�H� �12��x��9-\�	Ҫ-gK\8��԰lA��#�j�m��@P�"���Ƌ.<�q���Ƅ�fP�f��P�Vb7 �,�^�7��w,<P�L2�
Ǔ�l �3ծ���\�
��mn��x�)����ngCέ3Y+Z?�T,�źOTQ�`���Q�s� HKW�{&�Xr@�?-�_����1���U:�5��]��4�_���Q�g����C�WE�č���zJ�2�VD��¿	�F*�C���M^̆z��r�翰�n�ܢ.V/�9�����ͬ���Ք�bP�/e�Bn�=P��,9f�M�����J��!OٱtqzeN���fEFх�h<��)
c~��F˯��� eƕst��Ƨ�J5�U46&�2��9$rUywq�9�O���K�tq�􈯋��LZY7ĉ��6AD�FE+�~�{��#'p�~i�9
���<�r����2*����Y�	���(���+DF�1�5ʭ���y�d�M���nټ���y���B�������؅GZ��P��Z�)�-�YZ�V��#�S��;8pfv9���j����'?�n��������esk���bmn���٭�>���zKmi^�[��q��?x?��ݗ�G�?��!�k�ݘ&F��X��D�sG��i.�]7Ж�؛O�9���%/HG�K�Jy�e��g�d_�җ���OOZҞ�HW�zy����ҕW_e�e���[k�Yݻwo�L����B� �c8ީA����2��"�y^�ݰ���J���ؔ�\��[��gk*��[���?��nǝw�Y�Lu���u���L1:t,}��o�W]~Y��^�c�E�v��7���^��sy�ө�ix[_� ��~�a��f��^�yeurzs~��=�����r�<��=���i�/������#g����0D��4���>�)Y����#V�vTLPp�+5�X��)n����ЗE�Nc�qJ�։�QC�����ؠ��u-ְ�Tknǖ?�g�G9u؃b���'���)���b1�����N����؂B�ȩ^
�prα���'!��i�J�3ι���a���sA�ıs1�� �9y:�?�=}�Xp�:����B����s03<Y���u�'*����N�̯p�E�b���D}�V`+��8|	|�=((S0&@����	��e�� �[e�e����s�ǁH�n	"������ �hK�R��8X�h��";�v��^�Gp�嬈�H+�1q\���5�2ԉ\%l��4T4�6���a�އ��7Q�\3t�.|fP �b��ᝃ�������Nv*����BjYw��f����ԯ@lf(�G��� �l�����VN�{��\%q*nr+�I��X��"���suf,��g_�z���ԄH|'<ԡ�dF1.@.��`_��g�pnd�5�pv͓"	�ʥ���]\���ş'į/����+��ʢJ_ZC��#��Ӝ��|W��7��]8�� �
���fewEj��#")�P~�]��(�ΕIU6+� ��I��3�j�S>�1�\D���|�8�5��=���]a���p�|p����B��i;��^�6	�� "Uc�Q\��e�~^�vk��z�j�"]�-3]�����G{iFdm���wh
��H��8�J��<�F�vr�����X�1��j�j�I?H��|Dޫ(���%��� +�|�@BQG��4ơ�X��q����6������ѱ���2��Ӗ�v� �����R��)�I��p����2�h�O�ݫ�����#�8"9�����F����/�7�q.���ߚwu�e��뿖^�c�1����kSz�o8��7�Ⱦ�7�w��[k(�-�k ���]�Nw�u�ִ�#�m��������H�h�8��h���	b(�]��o���0��������@�����ց��g\��_�p��������Ke�w_�vl����KB1��o۶#���寚��q�����?���g5�}
�`�1U���	M��[~�8������Ǒ��7�o~�����׽.Dr.�r��l祗�n&ĉ����O�/����z:���tm޴ek���A8y=���M.�Mϸj7������4>;Yk�����\�����3���K��ᗱZm�Q�u�u|� Ëp�fЅ�Dj������P���;��"�.( ����r�&V�Z�� ��F����	��(�� O�!������A=Kibv�55�h��k�����s�E7�Sq� ����0���1�q�AΉa�ؘ���F���$ C��Po-�31���%�n�شL�������P�DL����'���T��l��މvL�N�C\K53��ʯ���}�xT�q��
�+�0�����b?9G�=� >��1���������_��#��yJH�&�c���/a�w¸y��1q���Ev�coY%���o�˶]�v�i5�-r2yi�]x��'�6� ���u������a�L��WO~˵�$�/pjc�g[W�4a`VG�'���qv�"3�\`���u Q6���!\��&�u����a6,�  Ǆ���Cۚ;=��)7��R�t�%�̡�6I�^�~�qf�
�t�q
��D��\�P,E�F�Iԃ@���W��^3N�!/G�I����6�0E�䦚,~8d=
\8"RWq�b�</�e��Nԏ��;A"B���ԗw35��V_����pE��ѹro�_���_�G��wˮދʕqh-Q-�B;�2�D����e)
R��bߢ<6���S�#�ʋQ��_Y�e�'�M��H@�� ˠ���f-����"ʃ����a�)���L� ���B�
}U"�4�9G��͕�.����c�<����&]���u�~�c��81]��X�"�S| o?G���[QɂB$�;���8����ĂKTNCC�5a\��;�Rp�y���Ӝj�5��qC�L
"
�X���k���E�
�H�d7���s.�ء��Ɖ0��:��d`gD�M�I�n��U �b���d���SzD�S�����ؘ�:��0ϭ8��ֹ�Bv]��A���c�8v%W-�cG�cg���Y6as��(avb>����&DZ��ʑ��R��8��i7f��#�ԯ�/��׿.]��;m�Z$b�E�Y��m_���!`�)��'��^��7���=�&� �eӆtɥ�\���.l� Q��'�%��ca�@0��`DDgIӹ�G�"bD��������~��~=�a��������K�8j~��W�>����W���/|���w���"��yئ����~t^r�8��]Pg+��F���VN��Y��|/\������DX ��jҬ���������N�Mco��q���ˮ��#��������pO�zKϺ�
 `!�y�`�w��T��^�����#Y\�	����bZ��PxUH8�V�󛯨��������R�Z�M?j��#�E�mE�b�gG���͚�M�3�9=L9��pt�,9`�g�V�3/Z;{�=c�n��]'�:;33�m�m���s��ߨ��9�K���X�X�gf�f���Μ�PGӵW_�8���Ԅ���-¹��l��1�0?��q�E[�l�i3�ˉ�����4s6��>�:}f]mb�6Zӆ۳�5kb.�4���!��Eo��jԲ�k�,��#' �.p�bc��3��q'�bߥ�nN�d'1_ �c��i��I�7������t��T�3����Q�'��-�\r1�Fiǩ��$D�3��a�B��;�0M�Q�O�/tM+��Cq�ݞ=�7r˂���0�`���Q��S兾*�S�ЏtN�=���߿?��B�e�S�6��n���z�A���Y�����l��X���}7� � �eK�}�"6.�+�x�#�G���R,�-��0}��$nj8�_��'��W�.#<�ˊ2�
ތ�
��%����X � ��X�m(�-j`Ύ���B��#g�!ꅷ��W�����o�ʬ�+"�z�"Ad�ߥwdl<%3�s�k�����ϋ�$U7WAѶ�Hn�S44�?"��+��wD�7�ߘ���X��i��Y/�8���Q�E�e?��#㢀"����A4cVui�S���kHƏ&��;�,[�z^�_��\l"����E�č��l/��4�D4I�2�}���D���U�� ^B�H"	"wS�btDf9��-�l|h�@6��Xe-�©q�8���kz�)�O�a���Qf���pe]h"]P��w:����F��B�e���N1��@�-؛��j
�5c���\'104�����h�z�����E���9��yX��H�p�a����3����M�Wr���8"��G��{�]}S��魓���|�#�?�O�����F����#��l3���Ɏ���8���b���s��K�A,ۦ���|]����k:�s�\O�M��~�ϲ�o�]�~�97�X �k��6������n�-��{��܋UYp�9d���مG�;6.�XL�;R����/�R�g����\X��q:
	r4�ٛ�e��p�׾u�b�e�d%�{��V�������L�a2��Ё�a����;��܌�^�Fp˲�8ѷg�q��[ $0
A�8l������L�%�pr��596�h��N���ytθw���mk����b�p2����)��y.�XE�\5!���4}Z[X�"��e�	��1ъ�7FH�⩲<w�q�9�Wpq���+و�\�Z����k�x&&oVf1V��pv̰ ,Xaٔh��ߺ/{�3����k�ȩ����A��=��C�-5��j�L�!�>�V�ؗ�fl�X16ɉ���l͐�3��x����lGz3��h�x�f�p�W���_}=ܭ����+��Ʀ�j�3��?`�ѕ�Q����\�!�Ԅ4J+��}�s�Q�˸N����:Fpt39_��X������� �>�1/aNgh.���A²7˷n����5��F��5����8#��u����zEڰ�0*Ŋ3�T��Ijn�Sj�]I�9�F�[�i8o�ǹ�jJ�l��1*�?v� ��Ke�e`���Nf�K_���D'͛�&��d���e>td9�;~K�f䮚0��ˈ�R����@"Nr�QT��,�ľ(1s|�)�6�	d��(̘ �RD�^��%(�_���3%���F�ㅿm�g\��������e�*N��u2��1�Ge�'<�������~*bUq��@´��M4�UE+Ő�X�`���쫂ة�f����r*¥
��
��UI�l�!���|���O�:Ve���ǣ�&T��+Y�G�Pr87q���_,��>E.�mG䪉@�5cVN�ؽ-�kb)�HB\�Mʈ�G�9��s��U��Ēy�bP�zg!���(�6N���N3�)³�^�J���˦VE��yay����a5����b�@u?�@�;iߩ��5-���ɞv��l��@�r�HQ8XD����dO��q{�Z�f����h�3���l���S�]��"��-\�3��b�h�\�]���S�ءwp��\0v�6���!B� �-��XpF9��¶Q6~|2k�j3�)GN�d{ߛ��*�&�ӟI���@z��7?{z,ۅ���_�b��Hc�����J�Fl堺 ���̅��C��,b+^����|.:ƾ"vc����G #��z׫�[]�1�r�N���EW��a$�.ڹbu��pّc�ᦜL���B����lӺ��A�|��ӳ�uc�Ȟ���>��A��1
��Y�f��l5��M����~�����C��U?���{0�u�����GL7=������Bn	��\W����L�D;�=[�/$������?阢oZ�۾�#z�((w�ŀ;�ѓstH=y���A�s]v��{�i���8&�r��;��e:h�E�$���D����#�3�[����i`� w/��w]��9�_�b^W�)�$�A�~�3~c����g���B�JwC �k�6f����p�T�r�:��=��?PY��)�w�Mi�ڭ�e;ͩ�E�g/(^�أ��.�d�b�C�YnlP���	aL|��p��I�h�#-�29<O�s%�&�J�ɡRl.!d�r��C��zJQ�ė�S|7\"L������B\��-s#u�ر�H�ч.�H�w�D�'͢W�N�M� �(u�7��5�?��Ƈ>K2O�F���~Y��j4�rW�9�!�b�!��`c2�Џ�T�(҇n&�*�����61J2~E���kk�ԥ�~��" ��f��	'&V����iXM�u�-�|��=�&�A!�~
"$d�r����N�p�^������L���W��+��"5a�F�_�����ͽ�Uax�#;�Ոk6[T���5~O�7�8\��Ƞ�Y�ъ�"i��`��  @ IDAT�T�3ИOU�h@�_ó�[ŋ�(�6�}��嗟E�ˤ��(F��y�q�Т����!�f��]�4~�~e�2O;���A{B�����k������>�T�**X�Y��wph�<n�U�Wq#���A��hA]��?+F��j���=y��֣ȓ��N�	��N�E���\<*"�xQ��%N�\	%��",��#��g�~QO�E��l @뿘��\�mԙ�D�.�Y,4g9�M��#�.�(���=?˽�, ��.��6��L�1"U����y⦏|zf1k�f����m���>.Lm���DD`�1^���i~x��������<�"s+����;B�����+�,�B�:+��֠7���y�2�P��zn�X��{�Ӟ7>�N��޼ysz�ސ�����o�X��3��/ٽ+{��GC�ϸ���t�M__/�~���x),"��A�2n��b"��!�U�V�u�<���V\x<A�:c��1���D;�ւE�Ep$CQ��W������Gǰb/O�X}�hY�>�Al��$�߱}'�@���~%�kͺ�A�p�l��]��C��^�~&���/Hw�{o>:6�m����c'�gk��ۜn�����t6Á�o>�H��{�h���pG��6��o0k��n8Mp���|����YD�^�B�K�̰�8�(l��*̋�P�흽�S(��������� ��js�f�Oy��\@L$d�qR�d��O��=��C�ŗlϞ�ܛ�?�.�� ,@d����.8|��ܕ0������ѱZOo�'���r� ~�.6=��w�G�	��]�\���UM��?�9��oߎ	X p�l��_0�*V��$��n�����b�b������R���9�"n{�_���O)f[���
ܸ^a5��IR�'G�іb3`���:B]@q��v�����9���������z��A�o	��cg�x�1G��<�����йrxǐ��"<�D�U��B-��f@&� n�qtO��gS���4߹.at�b84���)��`j����#�qÐ�X��S�@��퓺�ӱ��^��`�A���6[�2TwK��DV̅����֎~�X��;Ju�u�N�*怙����
��N��㿋�jM��̎��A>��6��9�b��Ypވ��r���IjѨ��l��ֈbʹ(��:Ţ*&�)c@]����9��u!K�U�E�U��o�c��6ILggTѣʌ���q�_4���E�����C��DƉ��;��ǣ>V�7�1�`8P��?�Ӑ�ٙԞ��+����S]$�D�����F�q��=�E�̳t�ĸW�Q^Y�2n�����u����7�2��,��,�;�g�(�6�0�9_��1�d��o,r���t�Y��!�W���&����!��B��K(V�έ��U���=s3�O
�?�S�ֺ9��a@9Rnd�҅~�#HX��p���2"�������Q�U6�P��qC�N����G��?0�m���C_��[��sN=e=,b�3c��n�t��yE~��a��`7��N1!��'� ��N�Iղ)� B<���}��rv�,���4�@���aa��ǰ��֒{
�bx����p�Ѝ�_�v��6.ѾID2r!��>���010����o�3�'�5�z��j�*{�5�B���B
#�O����wϣ윻�#�<�]�u'Ͼ�9�yڃ��fwO'���:a��.��:��y��WX�O���=�(�#���d{l_B,�ة�:{��=�{���8�;q�����"�_��gf;8�7������g]�C���K.�Dߕ��6�i=il��o=�\<��*̿t�j�ǳ.����>��C���<��4��/b�r��\��	�,�і�o{{��|��nL_������{܊C��S �m����Ԣ�M�-,@�@v<��b���{����j(ȣ��P��ک��7"΅��C�p���T>�u ��8ܵ���ϸ���.ϒe���~"y>���q�[Z�-�^c����v��g�!=~8�dW(w�	�e��#ںuk����ve��kk�v�U�A��G�FG�Æ������=��m�g�����9:`���V��"u{!��g�W��&f{{:G�����hPr��k��i��&��Xk����4���~[�PZE�v�Ru��gSsWW�"\i�΃*V�¹�����|�e�.���ޱ�"���*����#m����"͘D�X��3>6���[��0����+lP7��;��1=9�ɶ&�;)���a��\�ƉL%lc�=}�:Q��{���K�8�nB��ڏ�͐Y�΀{]�`��J�a�#�y�0,�n�@PI(� ��3��˦(%�P*��B,h&)W�.�`m�Z� �躿ʜ�. .�.�� >���h'0G
1! ��,\%��ɩ=%R%���W�)񈵛����y�x��H���q�f �r��>�#q��<^�Yz�U�:I�u��OpV������$��  �bWaF��S��;�w%�Vm;W}�ڈHb]c�����da�i�c��k����k��~|�W~����˯�;
�GY�3�0����X�y9W�U.\�D���+kS�Q/�TExĨʪ�\š'��Č��Q5B�3.�g�#/�Ѫ(\��:766�G� m�����/�E��cp�*63�@�h�Q��DQ�n[�e���1���X4Y0���fz��2��V���@C���R��)��Ǣ�Q^}���X�u��K�q"�#��31�N�+;r�wy� ���\,�Aԅ��Z�(W��k����ᣈ<zW{z;j�3K�7z�m'�$4�����=MCPg� ���$��)t[�.f����Aė��v��PK� �4�0�#Vc���9N���17�ٞ�QE3�T㮲�R6�b��/|1��_"�m[קk��:}���n4��H��;_X��gxj0�w#�>���.q/��"*a|���"7�c��)�8r�}��}�NBLۯ��wp��.���I=lPu�	�l��V�'?�w�艣��Ƥ�*V�/���r��T�����S�������}-�Ѕ�^�lڴ%c�vD-�1�@����z�o������9 J����LP:�91���������Q��`\��'c�Z�m�&���(������t�)�4�uB]�6�{��ى؛�a�;�'�.`^�zG�w�y�*�~tp"�o�{��m-��4?���1uAMBC���n�H2(FP�F��̡�=���������Q�O;����t��_8g,�E�oVҎ��v�&�8e?�s?��~ˋP�>����G����|px�2�����Њ�W����ֹ;�Ko}���W�Y�>{W��7^}Ž�lK�Ņ�~��sw'�T���o�ʯYB������۷�[2̱�������~�Ո�M*m¬~u�m��f�g5d��N���nOB��El��I����r@[�$��Z/���.ޝ�H��,"SHa��c~E-�@p���G$�V�Bs~Y_�7����[,�.$��s�V�OH tCe{DԶ��@*�E��ȶ#���e4żE�CSX���/u@sN�"�����A��a�QN�Z{+���Xa�b�%�c�<˲�P��i�� ��k���zc�:�kb�"R��'y��hM�-G�<�/7�QtC&ZYw������4�������q�(�^~7�э�"R�������cq+�Uy����(�U-~���i�˺��#����,?�P��Գ�c�~ыF!�ʻ�gY�h�:x��F���Q�D�_�.��0lf�*�z�Y�V�a�GI�G'R��Lc�˳�n+��w+@�=���D�,u�	�?���P������&囲H��H%o\�h����Wj[i#�m�48W`A�otJ��aqSn�&�$]���q4�Sm-ȸC�;��������p�U�E�h�;y��M�o�����o���ɉi8@\ʉ^����������MpKz�z��F�b���ZZ�Q�� LO�����i:��&N҇\1�f�N�lA�iyaZJ����иp4oV{���������b�����W1����PN�-�����0��2��>�/��H����ޞ6�/8�E��<��l�%�9HS�O�8�M��1�8���I�x�С����M7�d�,����
�z�!b�������}��8��今�Ɨ��Up���/�k"��~�D�]]��{��}���~	
��9Uu8m�v
�� �F���d;3�a��ڶ]WCԮ�������oCtӔm߾=M#�Ԇ��w}��u��o]6�AwPɶltj"s���Q�E�E��!�[����m]K���Sz��ޖ���M6x�ui)�L�X+�Xl�oG�C��xt�A�����>d�C$�VCd��p%Ga;��V���5�m��6�\�V��qEdOWom�qPL�zI�ޝ�r4�8Q=1���*���Ѩ��)�ʳa`���8�:z����� �̫�����1���ރAd�8;����h���oM�}�K�]�����O~"m���l����R��.�0���h���V�F���a�iͦ��6my�_s�����5g����y�P�������y���g ���y�)!u�#/T )���𧻓�d�g�!(�ˤ���5�]P~cPjvHQ�D-���)(�@� �&�8
��w��rjZ����~Qs򩭩-�Ch�C%y��J8��ǩGR2P�(�� B��>`���f�"sY���/U�'	���Z0���,p"l�e��ں�c��a
H�'��l@A�d( �A�b���v�M�HS��B����A��Ȅhe~QwA�+�Y=�O�& +�&�^OL�R,>��Wũ�_f^����>���_��_����?���������_�'���jۿ���b;]�m<����xU�m���_T>q�I�G5����֢z�4:/Y��e(T��J�
q�D�n�y�R[�*�ڞja�"�4�@F������m�D��[X�^F�$������|���cᢌ_��w�I�y�����>��_Ѽh��Df�X]N'�>�ul��p���<�FI�[�;�1�&.v��� �����y
ӻ/���l9s:��+^�1��495��oYWh.�઒��X�㞱0�A��R�����QU �U[85mA�`Kx�v�n�n��� [8�,��|<��Lx�O��A16���M�#{����+�3���$�zX��s��,�R��Ǐ|�Ex>�s�=��c�v�E�<�hڲukv�ӮO����za�n����+N/$���p���O�P�p�΃�s��˩B��8*֍�?�X��@��~��8m�6�}�5ث��K�6lN�X1W�F����y �q�� ����v1@?��c��G�i��B�k_`y�������S2�f��G�e%r����Y�R��ݞm��U�W/�hc��{q��#�W<��l�#�Opu�#D�	��d��<�0v�%o��8�Y�	�6��˾��b�O�6��s��W� s+�3�'��W7��\��o _�Q�W�X����Kd���p �(Z�Osl(��mO��Jͷ��/=��̊��x8��\8P\R���usx����h�ð%���0�q�=>����H5�[{��ږ��Il!vk(�Y�X;�6��,V6���QP���7NՀ����ʿ
�y���4��{�o���3�1M�_֘G�q+W�7��{��;/����xȮ�� "E&KL	f���y�a�L�]))��
"�X����8@���� >�|Ht�Q@Q�D�Z�v����~�<b�#F�D�`�pj�ҁX���(���| �(�<�������APG*lȻ��h~47j�$~(U���<��+T�ɺ�eH���D<�W.W"��h��ǲy��g�91�w6�L�V�g|觫£��[��W�׻JO�a�U|��w|�K�_>˰z�����0}�������<�����*�zVV����*(�F�Wm������hSᏬ�\q�-���b$�����ro"���w^}�8>������{�:ñ*j'��[�"�2�:x�	�6X_a;vp�E�]�9'(q3˜iji�I̎�';U9������p���$fP�"�ET�t�9��)��sB��tƇ0
�o�$�D$${�#�㑷y��d]���r�V�a���!�0��,�Sshg��X�w�I�)�4�.���������Q�~�S&�s��>�D��$=4�&�t>��;po3��l�?ۢ���3���Y ���%��X�xD�����8�����ap�#�R�c���.XN{>~8o�k��>8���_r�릴}���O�W�ޝq'?y�X�uˆt�}�Sw��9������7���3gF�āG�v`G��r������/#AcE[�rao�1 (�T�\=�w���]���a���A:s����@�h
�G�'�d�޸y��
㞜�ƪ�V�p��r�U�Lc\��(���mGT�����鸦�.l�5��.�"=pj>�|�P�,�8���֌���L��^��W����=\W2���[�\��aL#t,�Jr5�����w��ac���PI#����则&�f��໢Я.�y�7�*��kg�	�b��~�@�:��q��կ���>����bȔ����0#�{�+W�h�@g���'�S`�k��M���	hC6�a�pW�ua�i;K^��
��QK>��D�f&]}���9����/ޓ-�A��gX%Op���4e����u�\=5�-� C�e���ct��5�y{G;f���+]�^=+�Ƨ�fxc��z7�S��_�U�_ŭ���J�����G���@
��K�]q��3�8�a��� !�#�E'� ��h(���E��j�1�5��i�̨�����P�nx��&ʬ�n���Y�o��\W6D��0"WlzI�بpޗ�9���ܘ�}�T)��'�/e&�Y��«�|��>���}��x�{���E��\e����(_���:��ʿ�]���m�$�����ݘ���X~�GC�(���ק��B��nh�i�<�
U�OՇ��!]���*�Ti���y^�xy��|��y��W��yq��u�j�q)��(Nv���b�'�%�I�܌�#ʑA'2ʒ�џ_j����:l�IB"'\Gy�K�#��?Ɠ�AQ��B�V�ob�,���o�[H��X6�H,ږ_����_Ғ9G���Ǒ�P����&Mq�M�>�LNͥ5k7b�@����dz�K^���Y��a�65]�i7Y∺E����.D$���jT%�"ːc�2 E�o=AN��qr�Jm9��uB>:�=\����g���E-i�������� *�l���)+ih�����0�cz�]wiA:T�"��A���m�}o�%8�ܣ��})=����U;�7�0V~<9�F�"�lI�Q+�c��~�HK��p��?��}l:tP#�k ��8�>�Πǃ:X�-��ⷽ��3�sitr1�w�d~���t��.^���nDAĘ�[y�o�4�ڸ=[{��4�}w��xI�t������ �,�
3�~Ρs���fF�HB�$�i�d@���`�l� #�M2��`a�(��B`@��A0�i�fzz��s��s�~�S����?=xx����{o�:u�ԩS�NU�o�?=uo:q�����ل)�h��M0ltv8����ۼh�]O�x���w��v�� k��1�A_��>�3V�9�׋x@��T��F)�����T��G,�������܄]B�Mm]����T�H=O;�%�t�v:r�8R��1X��p�����T=���h*��?�,
Џ��J:x��Fa���9�I�kX+_"ONyVJ�vz�����Z�J	Ӓ��h���d�M/��qx�ِӟu�?���*`��h>܉���n���N����?���fq�y}�x����Ns�<�c��W���CF�]�!ա�p���t��Y�A�<r7��@$@.IhL&��ė@��V`�+�@!�t�����5����y�bl��(ヰ>��"'6.�,������R���t�L�K�x��ՆE�`j����<O �T^?�$qF��ͱ,�E���t�IN(-����kT2����M�|˞��~e������	�ڍ�6��q�n�Żm��{��n�-0FQ^���:ҘO 8��lo��������Ƿ����LZ/{��~g6�Z�����W��F�>��C_�E��D���aٕ����k�|b��k��y� ����Mq}v������$���l�-��t��!!�IB�Q�X�\�"���9ۜfa�%�܍202W̫��2[���sxhy�ǡ�.�v0;n���A��-����q����d!�h㻌	�`�������w����1�ZG�`���wBq����fJ�ap�m����8���I�e{(ś_^�9��{࣫���bE����'��E��UƂ�6�T��d��BM	Tl�tz��%����u<�ޚ# �P����4F��Q7�k��5�g�8Ϡ�2P�pC��rO��w������~՗q:�P����k>�w+-����1�8S���/A���˗�[o=�ti:$�Yڮ],%�+^��� ���m��짨Kf�����k����h@��I6���h���q�h\I�+,N���U+�k�h�l�����c5� ���ˮ2�!�Y�DJ;��`LL��K揙�(\���c�J�2�����j����k0���4�M3�#����Et}���}�!\B�g�m���q_}�p�^�J�C^E�"/?�ـDhP������ �[W�:�%>JD���Q�t}�O�^��/L?���O��^��O���5r��&>�����ݸ�>�4s�#�,$�U��z1�:��t���t��0�xϽ���{����8[�n�]z�l���>�>���ٗi��O���5>}q�f� t��-���=�8����DA7�UEW����7FzN�H��,lr�G��|?㵝iKXy��m|�Jx;}�Y��ӿv���γ����۸��=q�8x��������oM'K%�{p°
ѝ��� ���P'�s���Vrl�O�QmH��.�'r)q���m9ok��%���?4����xbe|kȔ�$�F���7%Ĥݤ�ͯ��.�5`�T�8~r�����xF�#��r�Q%����v�>r3QJV��i�aʉ������_җ��w���V�|�������Ѹ���?�lA	+e�wd��>/��<~̦y/����]\;N��Y�l��������O׿��z�Ky�7~>�y����哸[~~���a�r��|��T���4�����`n|�-�pe�
?c�F&M�'8��<�a00.�X�C#N��e#��lU�Hz`r�_�x�� S��ɉ�r	s�ƥ�F�=�%���e��K�vT��*q��:�-��,GI?���^&Z�[���V�|HP�G�'5zF��ް.=��N��됆uDח�/���-o�.a'�������g�pPw
�I9�S�UJ�ʁ��N��Ǩ���3�L�:OD ��ŷ��L˺x갲��2�Τ}�r�x:'#c���J�]�E����a�ҳ���Oߏ^�B���Vz�K��/��(C<t�~�'}f�������H�UZ�V=B#yr�$�^���+��𳏁e���'n�?aظ�K�h��+}���G�zf�ϑ���#G�U��+o�?���[�K�����O�o��oI���Q�߬ǎc�혶`��F��@�4W�x�'�X ����A���W�  ��v�q�B5̔1{�\Ry��
׎�atay�^>w���z�~�+>7zd�Nݰo��Nʡ��m�mh�~An���D�Y�SLx9�Dw 9�/��t�<�ɦ�=�X��p�Hg����_��f���ק�|���y��l�pR�v/!�D��a�:Mqe��º���c����?�������OU#&Ш"x�;��i��|}�^al8����_���I�&������~�z�ߛ:\y#>{���Řt�fL�u�g��1��AwY��Up&�3��a����޴>u{ӖrJ�Y�K~��f���-p�K�|p���sy͟�O���,%v�¦�����$�e ?�rt ��wC3�å8\���O��?��J$�u�g��wĊ<"����@�y��`dB�$l:������cދZ),�	��~�������PmxC�s�"v�Q�x�� �����3��tz����de�Q/�����R�X�V��������2/�Q�|û����_�S�D� �4/�J\Ӷ�*u�����rz ��=�����/���z��zE���{�4ჟu6,�̋�MX<�T
��U�7a�|QN�-�������M�ν��}xC�Mz��[~�AƦ�N`�-��ɸɅvYq�]T	���2�yqB)���c�-���Z�'�d6<ͦ����;�0 �[V�[����j�`�ڐ]%��a�1"g��c2 �(,��E�>�P���#=���e�t����^S>g�(��)��k��	_FL�d�X�.�5��ڭ�,�=v���O=�n{���1$�������r��g	)���ޓF���d�k��S��9�O�a�� l��r����-)1�5!��+o��(>���䩿���0�h�E���aUgh��<ԛ��q���= TQ
tuv)��o�A:�-_�%_T���{��a���/���c�q)&R'ȧO?��N?u&�z��O��(���Eߩ��d�KL�,Q#�٨Y�.#{�[��E��=N`y�y�mP����Ҏ|���� ö����D�>���셨d��q�ᒰtuq�KS�9D�>�F)�]o��8�k㜂���x�<��<< �a��^���_�><0���j����D�'9x"����c�	ݤ׼�v�a��L�w�H�0s��]N��N����n���c��c��%J����)qA� ��#�i��4sl�x`^lŎ�Na4t(=��������ӡbhcm'�C�}%�G�0�@�F�(���R��A�܍��ELWLOc�#L��,W�!7��Lp=zy�^��гҳ�j)lrZ��P��o�v��F:��ܟ_X�R�Z}��[����0����A���������"��2�/j��@�y~��8�h4��_�����.�ZIC1x�ϯ���S���ް��%^ɫ�6�%��'&c8�!b`��Q��ĭ�3V:�2�k1m�J�2ێ�A7�$] lMsb��',L�Ȇg8��Fg�.��������[�"e4�x!LTr��%�̓a��#߬G�3����,Ac���'r�A���vK�]�;�3���nuiNpM�MFX)�<ͮq�u_<y6��5��l�7Q�۴ů<�~��o���gD�^�v����m6������x{�4�f~7�o�7_�u%N<K��m�9&�M������17��w׻���=~~v�l��A�'s���TDN�p
:�)U�=޾]bOe}k5N1�#ERB�4�.҂�G�m'�uR*�#zH�`@b��-�7�AJ'dN�{q�u<�h����#��/�b[���$囟��J��C���6@���9���`,o���vr�2�u�k��
����clW]Z�ν�k���'�����C����j�+=<�͉�X`���Q�M?g�0T��ŗ��j��l�"���r�@��uv����h�v�5��C�j{)��c��i�{1 �h���縉��]���M���ә�������xA���H��=q'��B�7�Wo�_?��Cq��Vŏ;V8|�~�`�dL��=�]�M����]Ƶq!al�Z�|v�Ɉ"�����zcJ����s��^��'F*�[�O���"��<�����+�q�[Hl/s��*3�& ��+0QPF�V{��W1�}�����I��ɟ���~W9��Q{`)Oqv'fq�(E���z��r���G��3?1]��f'�m�[~Afct�ɓn��{3N��3�$�J��R�)H�q�k��q������髋ՓO^��>�����~v	ǁ'��.\Z�W�a�ɼWq����`p��no-Է�<��|'����o�Ø�X�#��:�����V�I���Y�;���PZ��^\�>��U�z%��O����2�%�Q�$� c�p��G��x7H� 1�2R���a�V�߁D��}��v��q����(��8�0��~��{��u��D,�䅅��c �Qf�8f��)��T�4D�������̈́э��� !����C&�\�+�����}׳�"�������9,���U���1��u����3HX.ؘ���y�C��p]�˯��cqV��L��ϊ#Ƿ+jÝ�p�� �e�0�P�vMQ&n��&n��QFI�<�_y��v+辡|�E��#r)�<MO�E����E=y�v����p��%P��{�?�uC��k�'�z�v���Q��^� (S+ߦ}�h�S[vM��g��J����kG���7�_x��/�H�^�jS��CQ�BO1I*���X��%0�򑸲<�������U!��$E2 N�.�dnX�Z�h3d;N�����a!��ծ̘i�{�P��`�x���5��G�0�*―Cql�u"O��`�vT<��˥�����f��g�9�����n��B��ɮm���vW5��d���1�8�vǇO?]iix�ɩ�׳é��<����6`$71"���^K��'	����no*`w˞�,c�l�;�
�d���j�H�v�@�����
ǌv����D(53�C�u=�=HO&1K�\�/i�2������+K�����P�^�-��C��4O�I�[n=)�R&a�°W�Ȅ�'����iQ�>���o�U��Ӣ��~�|�5��a��X�f�3QO�[O�~�w�Ʊ������_&�����ʹig�w���v��Zc�~�ؖb+�O���Ö�l݃�����O>^�_>��bU?�wS��;���!Ҷ��0��R�uHr� 6��Cm�gЋn�xm�y��2�P:|��ң�g8R�m�L�\��,%��i�`i7�L�x1�����%�<�H��2J�W�"�N6jL��ˁi]MӇ8���3u�p�&ȁ:w�j5
����c��gv�_�Z���Ɓ飏}�>y�0��c_	�������dZ�Q��6? -�O'OݎD	��c�Tׯ����I����ܑ��j�����i�ׯ�c�Op���n5R4���-#�1?��HD�5���9���)-?�BP̸��{O��,�}_��W�?�wI�����%�����.�ӛ�c �g�t�U��]�œ��r`� �ͣ�h^I�&�++�1��L��`���o���A@0��r�ޮx7��M��	B�q'�<�������~���3�f����.��ہ�w	�8�OO£6V�Eh��4��
�F��gD�'2��9\�Sy����s$}�wis�`�'ʷϋ�/tM�K�Aa����>�������[�F-�����T@��Y�V�mwQ~�#]+�<���7K�y��oJ4Z�k�>���R��lFV��9���fN�Tw�B�=;⹥�d�c�Y�״��\%O�5����ɤ:���R�[r2[O<��8�V�'?%���~˴�y��z-��Qf\�aYJF\Q�Lq4|���5���a�.Z�����W��������1�<�2Ud^���vܴwe�܎��Q�݂iRf]�����*��^!{�z��=*�&���KmO��߹��+^W7�����`/���4�F�j�C�Я�+�m��q��gfi�z:�؇�`6܆�r��-T�G"�]TJq�,	W%o��w�U��S�7q{��oX[����s�ݺ�~��Xk2t�`�3�Q�i���g��$��7��[ҏ��K��i�M��o��d�� �z��=�����د��/�O{�?�y^O�}ϟ�G������g}�g��������XH�F�I���T3��������B�0��0108�����0���
?�Z��+�������<:}s����;�Z�ߘs�Ka�v���� �1	�C5~�#�#.���E"�uؒ�h$� �`
��t�-.���>������^N�;���q*q|r_u���������8J�M����̙3i����u������ى]Gؗ�U�8��?���K���tǋ�O=�P�����;��:|@�� O��;�����N��}?��&�^��b���8hk����*�_�ml:�J	\kX�]W�K��m����j���)>廤i�Wⴟ%�f����NW�{��v1�c(	��:|K���z�F¦=E	%{�C�tpV��¢�a��W��-�p0����z!9 ����#�H������V�Sq)���z;x�~`cJ<����6g]��Ք�]�g:��4��-�TˬvU���"���EĠ�q�m��8�(@7H$�~N�p�
�OjɛE�6ѫ仫�aYv�էb8���̥r�a��+M��!!%��4,�������W�����.w�FZO^��P֞.��RG�<��p��=W��c
����J#|�HK--�}�&�n��å>�@�^M�����\~w��zR�(�����#GH�C�h=��M��L�S�͔�Ӊ1��ٔ/9��p�A�r˶��+o�=f &�e{�-�\Q~���$��g������%^~�L��E$��AO[qm��������&����M�N�0:�U��^Fo�;԰mrxj�����jmqy�lP�1���=�
��ؒ���i���w��t���ϭ%��~1�*�c���{1�i�u�-����i�,/.��G�ö�ҍ�J7�E�_'�e���0�1
I�PÓ��b���H�Q�ŞRV��`Bl��nx��p�|���N��ު>{�:���ƪN�1ʸ�j2-3�V��D1y��=�~:=y�R,���F��$���l��� ]�����v�~�"��~j��� Z,W �S������v�
�LK�s"�ĦPu�VNH+HYV��j�b��-�af�+O��Ǧ�W��^�4^/m�WK������	$��3�o�M"�`}��R�4j��r>15�$�SX2L}THf�J�D?�f�c�(�#�!h$���x�O�Mի\<�).��W?���\�.�W�߷����_����|�ק���#�����t��᣷xY���������_<W��������;���~.������G��U�9��-����?��T��c;��	�$�r����U0�܄��w�a!�h_���]�p-�<����D�/*n��V{�&u��|�G[�S|A>�8�t�܍dٟW��� D?�=�t�=i�P
�i`�b��tV��^_�K뗟H_�O�>fg헟��KDC܋�͵$'�z���TG':��wd����Χ}�kӿ�Խ�q8�kc�Z��{�����ϯF��o�o����W�<}˿����1��x��=�������~B:5�ҋ�ܖ��������4v����Sz��#�pyC܉��;88�چ�|d��e0��(	G��P�9v�-�{��/i�aſ���2^ɯ�������V�ѿ��$�
VQ���>Zq(2� 5�H�f��6�$`+����b�F�s9cbϾw�kM �X���Zd5��`�%V2T���0%K80ԓ!�N�R�g��(H*/y�L�*�E�3���F#�	f<#�d�x�ѧ��P"�����hٛW�p�`ؾEȶ��ރ������z�X>f���\<h�v��<��-���j�.��U[Us@� F����]�J%�JVR Pq~r=�l��������"����|�ɪ[@+M�/"���{�2��Qd��y�/��&`O�����}'j�]�e<ѿA�_sY��.��{�u?�x�r���4F��v\ûm&D���M},OW��x���:�]:9ļ�6s��A{$'i���JQ��:Nm1oUsܤ��c�025E�k�����A�!�
8o���7�s��u�~ ��J�t�����N�.f�����o�1Y���J��̽g��|2A0C!3�U�B�0)&��$˭/$z���,:Hl�Ȁy��[o�֑Vh�x��� B��ݯ>.�Eg�r<Ad��ُ��:��NX�R�<3F�T����獮|�}�X��/<34�fb  @ IDAT�Qf�KJ��0}�ux0�w�zAOjk���3!ʻrikHHF����ŧ�vA���j�m�������ܠ�Q�Z���b�x)Ps�UFW���	J��^zJ��6��G䳃0��`���D���HN\H�1��>�dz����X����������'Ƨ�T���� sAo�=w�_?�`���{ҷ~���H'}ҧ~r�8����E��C��O�� @��ڼb[�m����ז��\۲��Hܙ��Ƨ��#~��� ��,VƁ���S�G3��g��V�4��	�ĉ�옍^¿���o%���8_"�K�	p�]�Z]I�1�x5Fc�1�Ͱ�붥cc�����谒̄�봨N_�_� n/I��{�~�~6=��ǪO��פo���:yr8}�7}]����k�?�������������7��H�$v����/�<+�_�~��=��"��i�+�8~e�mR`C|
�%H�v��w]��_�&��a%N	/�P�ƿY��U��n@|T�D<��yh�:��Og��N`( ��AV����ݺ�Gq�̅��4*9aqaLO��*�!�{���0[�TX����� (:���Ʒ��3��Hn<B#���	�:�1�,����OR�U;�in�\5�5�		W���v���7o,\�\�����Y]�:`���ڜ�`�{?z	�O'�f�!~��a�Ë��$��R�1�*�j(���z1s�n#"���EZO^õ���H�%j�8Q^Nd���{���4dKc����|�y?�~M�y/���}|ӧ�򣌒�����Ets��EM�M}��zHG�s���� mT���>�%���sC}sXS'���u���]��N��ؼ�ݴ�մ�)7ψ졮h��SD�ԕJ�����ul�0=�L�ս�,`�z8&<�]�ўq$>s0���y	���H7��kiV�܋�tǡ�x&gKt�¬�B��Ih��'0'Q6��Tm�u�,������H��
	,��bt�q���K�])p݇U$C�/��v6؎�H�a�H>���)��؍	j4���R���*�vh�8շ�<U=|���º��VP���H���*떟���v	e���
~i?�ŭ>m0�M���MtC�|�HS:8,5Sƞ/zMs���P�]��Zv��.����.��!��2�dl�P�uN@M;T�gV�|��;�!�F*X!
S\E3�m��dm�G�H��p݃b�R����j���������2���yD�%P=%|$B�
�x�Q�_p��[Oނ�p��w��T��w�/��/Ahޝzp����v�b8���o/K��;�X���ru��o�<~��⾗��^8}�Z�Q<r�}�a�{��ә��	�A*0�t���;^pou�w�ۜVD��ݢM�_�~.�uΠA1��FE�����Q�.��E��e��xD��A���x���l���1��7ȩ��#C؅�NV\���u�t���ۛ�m��Ó�*\V���ru��H��u��R�/?������?U��8v���}_���������{��G��w�=��C����;����֛��?{�l��?��꫿���Y���̭��Gn����C"��N�{�H���vqqm��8�'pp�J��=K�̣�)���[q����]�����cU�7�V�[f(�����U���\�)N�Ox�+ӿ>��c�IeB��;�M�d�cr� F�%�6v5VA�����O�F�4O$6������5LO��W"L���8}Jĩ_I��Q�i��掦��|���)�k(~W������Y�������b5<̀�*���ܐ�;:Q}���4�D�	����Gs";�=LJ�pZ�]L��q�,Tؐn9Zx��ް�;Ǳ�f���:��#M�[����/���&�������P~7��K7ҕ-�܇�Xߦ���~�4ݜ�GP�Ex3����u�Q��J�v^Q~0��:���nv%}�Y��~N��<!u���r>b���A�$��q�N�C(�2�9������έW��q�s�����'Ͱ:�l{22��>�OB#<V�~4~칱�L\�l�+_�9���vZd��	mp{0�2BQ�e�(�;x ���w�D	���P�o�ճa!浌�\\�;6�cxt5��2�?�H�ڏPfqm�;<�]\���K/�U�}�YFI��!l��:�t����SHm�L(s&�q�$(�Z�V��}�g��5~�ɰ� `�A#dOv��n���'˴��1���	�㡑���'W�R}ÿ����w�U��w�	�l�|{e���'��t �����:; ��6?�6F�CX?S�,�G�U�r�_F�~G�z݋�1���t��{��x�h}��I$yZ��H�~ן"͸����r��x��=w�ˇ�����yYz�O���OߕN���t��>x��v����cui�'}�}_���;�Z���5��D����i�q �>��Si��z�����җ�"y����SW�����?��C������k�n�����,�]^#�#?�4X}:��!��E�5g{�;��1���"�gkli~���z��k�+�~񗫩���ǯ,��{_����ӧӧ���&�Q�Cڌ��9Ͱ==�o���@�:8�n���Υo���
�H�"��ZD�&&m�x�����,$\2���n��>?K8�0��5��}��u_K�V>��̤����7a��J�G����g�q0ͲrZ��$��"Y�s��Þ�DU���z0D!��D_0�[�L�_}d��������T�ɦ�>
򕧝���]Hd���#�H�`b��t�9XՒ�|���/�DfM��m;�C&cd�AnZ�����%�{��g~��4����R�h3ԫ�PrC2���s�;��0����tX�B��Q"BEb�ꎌ�ؚζ����ͼi\�
�2�7]D"N	��wq%����!��Վ�K��bb	_<J:� ��#�7�����Qd�.�cv3�;Wϗ�7�Ś85U� K��+�����<�-!'W`�d@tK���PR��xy��(��g$�Y��gS� Vd3��K\ͧ�j7}�X���Ή���w�O���S��]�1�9�/�Q��XFٙ�"�rqӉ#�2.2"*c�H�m2_��+a1/��Щ#�!y8�+@���nx��&�k��Q,��`��20���,׉§nE]i�J��'����{�1o�4j̎=d�ar<�̽_wV�l%q��)N�a��+KV�di�[ot��s�Hά�����O�r�Xd�Z�"֋n%M7������������� �"b�cv��[PY2l	 ���6�&��`�2�P�����j���4��@��%���9�7Νl�J����gQ>[x���I��P�;@�R�����ǂ`@~9(a���%W�D��}��x�Y�O����/�`W;r<���~�/�o�:il����i��Xϝݹp�Ғ���C�	�Y?�s?�x`���B�������w�]͠�����Kl�a�|��S�5���t�ܹ��NA���ĉA��7M��&*x2�#����k��f����k��{)▟�4�ޔ���8�c��L�7�5�m�����f��ˎ��sq���i}	�����4@g:����W�p�d::5�^�i��~�W�'"��V�ӠOݙ/_�Ɔ1^��f;X��+�U싍=�6�ҕ�w�:�YZ��7R�-�����\g"œ�ls`b�f1�!� h,��XȀ�e��W���A�����MP�Q��Գ����_��^\�+�l���6{���`�K����k� .G\Y���*�;��I��)5i�e� ���Z�G��m�O�h9~�O� �/�3i@�ӘO��|o\�k		��R���G�&����Dw�ʼ�	�\	.���p�@�@� �}����qj@ HU�gsH%�cV����2?�[���,GP�ʔF7�$2�W�aL��!��Ǒ�E�'��sCԢ��'�=�w�q,�hd���V ��x-~��9}�3�ʕb��n������s�g��[�g��ʓh�I�K�Ԯ_���v����>�����+��[�U�BIo��^"�,���E�&n��Y\'b�1#�~�v��gI*Z��Hc@���L��z��i��f^]\���l�+�dk�\�pzYD���8�C1�������Á}n���v|oc�Y]�ʐt��Q�e36�zӶ�Qᨵm�� ��l��.��P8H2"Hoj���c�܇�ǹt�bg����qwF!��`�ԓ������_�����[�4��X173��I�Ɓj�#�\}QMs�|���W��Ɯi��V���5VAÓ��w��h��t}�o��Z�6������n��(d�j�5�n>���PO�ݶ��(�A v)�R��U��&��R�����k_4~�sU�q�i;7��X��8���l�djqQ�B��k\=yF3���r����n�5�Y��	O�2���_��W���-d�����l�;?2��{�O���O��<u{��;�L/8uk����+�T���ꉫ�p`%ۡ����Zu�hf������cO=U=��r~�����+e�RC��F�lU�㴭�!H�mnn\�~+�]G��F�;2"�~����t���G��Q"G7l���8�O{A�mp�t��R�FR֋�=�[�1���D�����c�>қ�:sh�Q���0C�3�Q�mv�*N�9��#U=}�Szy�Ǽ�2�2Aȁ	,}��H`ޯ��8��H�Q��5L��$46P��8T�������7�����������#�-a%��g	o��{����Jz�}��ҡ͠+�H����A��>{��p`0��������
�$$.���CU/��`@� �U��O*b�^�j1�GqA<9A!� �D��z�|x��x\PO�A���c�t����m�q����(�<p����rz0�e�9/�1>��/Yx��(O)�7�GVK�f`,9��>ef�_����?�{E�ALspr �D��`��^$%9�F��*�Z��AI��^�1�N���`��o�n\���.�����뿧����N�k��s8&�?����=���cT����|�7?M��(�Q�T-1N�+�s��\���[����x�|� ��SD!����o$3���ϐ�K#���"q�h��������rќh�*�h���+�js��&;K��"���N4���x��&�� �v�B(k��&��6�q��ɒA �hMoq��.��x�@N����7 =�-������4��!8���{�rh���aЫ�+�2+ׯ_�W4ĭ�؎��Vue�RX��P���Ə3���'�\���̑P$�C�;���q.�\���b����
�]�+���,��J�,��>��ښ�*]��m�P'j����By2~ů��1��v�O��y&�����dk��P:�l��&�v")��iצ�bց�/"!P��O�uN_� RG�j#G	A�ʥ����Q)�iq9�����DJ}�i��,�S�p�A�a��q��P���3Ht�����W:��O}ݧ���a��b���$�l�a��h}4w��y���v�}�Eu?���Q�x�/���S�X���~=u�>�����'�=GO��2���ٙz��x:y������x��pQ/��A���af*@oF{��h����>���\�D�_8����+ dB'&>��2���?�������f,�!.�lVיFlC�L�Ͼ7M`��ճu5|�B [��Zq)pz�ܕ��)Sq��cOV������g�T���:�:L����;C�10<F?0�1�������_��aJask[b�ig�B^�6���K�\y
im��@��k��G	ξ�|V�ƣ��^�����G
k������c����z���Hy(��酅�[u����Ct[���-U�J[\l��V8k�0�;ѻ�/�� W��`Ȇ�����IpY�[{�`���@��#(# ?�Mj��0��ci�����O����?a�;���R��� m���?4���59�0r�9v	���xK��N�1D���+��>�YH����3��A.��#l�m�)�IL, ���1�
e��q��Oxwqϗ�<s�]�HV<�<��j��0�7���o�ߎ�~oE�����/�'��<�	�J��ԟ�]Ԑ��o��$t`���`~���z�c��dk��Β���~3V
��u��Űn�t�-�1�G����[Y�eu�a�˗��q�]����j�:��8L w:)O&�-D��C��������J��2�;�Y��l(@M7�µ�Az��!$M�8��']I�1ڐ�:��4�����a�_Y�Sjʼ�L�00l�I �T��=��N3�U$n�i�[o��{�w������5�x�&:r�v���e�QL}fa�^��z�xك�P>�cNf�����d^O��,x�c��&�����,�u�Mo&�k�?��x!���H��X�2�ld�Q�hz�Ϭ(��H+K�qL�����(��Օeސҡ;�B��$��Q͢����H�� ce!�Yi�AA��j+�7EZ�>����,6H��i�36�HtW���Z�Gy)������m�݁A�%�|��3��$�"��r�J��J	����ܕff�U/���t��0�\L��O������߾�ߤS/{54W�u��	�Օ����t�ή`4t3���y��YD:�T��a���b!H#�7�/\ng������:� ��8�K��0����?%�ߎ��SW�������'�T[/O����/����c��?��wԧN����j,��CX�>7��!ȥjuk"�`E��G��n���!�����Źt��k殝�wP���MO:3�Pos��$&j����a�W�a�z�J�3���x�k�=R�O4�:M�0=n#�]�fx^43��vm`���k��ݴ>K��
�ߊ[�/O�]ۿ��N_��̯�߻�z,��v�(�S����ݛg����
%/W� |��AD��b�y�f�"`F|��zJ��%�3�!���� yw�)���T�ȧ� ��O\�L��$���d�-P��R�d'{g�>x_��A%;�tS�M	G	�'��|�+��pB�P� ��2YK�,9Ʃn�ނ�s�zLƎ��10��S�9�X���%2a�ˆ@Y+[&���:����o�����f�n�	rb����+S�S"hY���]W���7̿VX�K�k�J���=I��M�>�qV,ҕx������vI�࠾V޾�|��y��X�N��p�_�`W�v��M���^�|���셑�#Y��S�E��$��b��¿D�1��h9�y���ݭ_N�=K _T˶�2҈^���'-Ð�J���q����x�IV�=��aI*l�=��ȹ�R)��}�@IX��*\[7���h�n)�+�E�
��l�	�#*�����g'Ψv�ȞU�ĚB�ku�XH��G۸�	n~��C(ieC��tg�_�U?������a�$�m��?��Ƨ�#���~yq]�)��XC���
u�ߴY�ib,_��?/e��'��|����a ��5~�k�bC 7��|�(����X'��T�c�ΕH���gH��_�)j ����#l���Z��xuH��&u8F��)u�6�w���(<�����Uʰ��W��6.B�B���9/G�g*�$�W��'�����A�]�z��ƾ�����]�mo|Sz�G����?���E�3�p��ZJ�[鮻�L/y�}�C�z�g}Nz��H�<Oc����|��eL9V��as�I�2�_��������i���sRS�i�6�����p&w�V+��a8\Ta_2��]<��G!�;���Ȕ��I�[0|En�\���V������YX���U�4��P�{���tx�Tz��|J������;ҏ������צ�O�5NO]٩���G���{�<F(�u"������_���C��ix�~�������o�����/T��u_ɾ�RH�ZU��K��C�zM�\Φ�뫾"}�������ҏ�¯�y��Ƴ6���%�|=?���3>��&������h|�g���o#2n����0�4��*�f�_\	�o���|����R��ǪB�B�,�N��|L%ьglVC"݂3��ͥLHLL�����]�md�?&7�3H�bq'�z�k�û�g�&^@���Y<��%M��IYF�I�'�qAj`����c#��d�T�����F!l�=�!�y=`BK<�ܳ�!��Rl�������@1���m�fK@#
4a���+�G��)~{��i���v�� [�&b]Ɂ|�3�3�~>�k"�}��o��y4-��]�F>��d�[��K%�n�2�\��1&_E�n,��<3�����ėf��Ho:���������w���WZ��c\]�Ə�9��[F�s�S~+����iӂ���`���z	f��=W�#)E�����*�XY^��?�jC>o^��m(��Y�D�0���	�|r�Nl��U�\H�����2�^�������/z�Q�8�P����&��I-&_OpWl�y_Tg0T���X�@Q[	���Z}u��M���Oظ�Noz�/I/\�瞺��K5=2Ω'$\��Њ��8��2����;z�h��(��.���yd|�hx�,`�6�X��z6���pk��p-�`�%��0@с���}@Ԡ�F&�A��B*Rw�� ��ð�����<͍�)ƊW�8)�6�'���ކykY<,�-Su2���b|�)?ǟc����4u���([�G֑���q����Ρ�0\}�?�\�ez���Z���"��0:��K_R{2�3��K3sh�U���xGz���'O�-#�z�?��?�H��j��miQW��G��W�\�b��1��5pha�I	�u��;���6wű�Ʊ䦍 t�\]E�e�ѶҾ�L�W����1��o�����p^�������#Ov��P����[��<�~�����}]u��X���N����G���o������zx�(v��H�OC_k4��ߜ~񭿎$o�~9����0Z2p����V3C�t'��|wz��������^��WV��wF�^v�x࿛�b�[m���	�dx��������������_�7k������y��M�|��b)�,�T��o�����H� ��ѐ����S'�%M,��L�`��eb�y�`����Q��smWD��RBLp�i[y�HxA�!�:���,��nF~y�����[�|�&H3	0	Q\aI���Qi��B5���f�6��󔂈$�~�ሄ��'�*�hR�d��hk~*��~�W7���M+��B��U��۪�e��ȨWDgd�z6-�����ZF�Ⱥ5����D�)Z�&������~�r!nȓJ�!a�!Nuё�XS��gM�:9�x�5~r��Ԟ�p�m?��km�@ԝ���z�z�42�����<Mb�r<<����
	z��/|J9�H� r�/]BO�r�9rS>5��u�#��٦�8�|�ڌ��5��H)؏��Ig��^Z���V�����|)�/Z�?0���B	�)�C�����{���%u9��� ���cL�0Hċ[ ��ȟ��9YQ�Cg�ӣ�OkL.��J��>���1
����ox��
ʃl�[�G 5Ig�.�s�f��=�z��$,jb�oi���h1���)��D��+i�,L�~�,s{ׂ���3v��'�m'Z���i?6mÏW`�3���
W��.s����7�1�
_e�d��%�`�,�M2���1�����7�i@��>F���Tf`0=!�v�͘�9THBr�-(���[�cMXs��29z�
�3�ϼ�/v��:l0��nx`nt��e�)��������;�Ip�v���^��P���rkTɏ������9c6��>�VǗ��^�$�$���������ׇ��^����`߉�#E�����Xf��j��}���'\1�	ÄzƁip�F����� n^	n�R�M!���y���������ŉ:������ �ٻ�h&��������ߍI��_����?�X�L_�e��A
���x��R��ߝ����ůz]��G����{���c����x(��_~�%G�a���Z��;��7T���L}Sz�}��ƪ���T�F�������
�i��4�jjB�G�I�vǴ�9=Z���]@n��o����q�yf
���u7��U��gyo�i���v�Jx)ߝ�fʐ���ΕFl��}�!J�%,�3�q:9g�0��"9�9���3�Z/E�r�w��<�����o
ҎU���3��	f�ݦ�r���Z7�b�&���$B˔,d|��In���li�Ap��� �4[��a��K4��u���K�A�gf���	ox�Di��~�+��Y£}մ3���Z�b0��m�v�ޣ��Z��K��|��)�Q~;]	�=O���Y�4r�Olt.�����C'v+@0�I�i�d�D�1�-���Ϩn�gh|�S��E���//��y�r��ބŧqK��I[`�7m+ʈ�g��pC����v������4�e�L������C�T�^\D�ہ��ڭ���/2mp#�@��N���ΐlO�m��X&r��Q0ܑW�ǧ��}�x0O!dܷxǂL�
�y<ʐ�]o03L��qT����e�l�0-a���=��%�f�bs�@�?~����TO]�����d��Ĉ�B�QJo\jɛ�֋��w��5�D52r ?ЇP�nP�4��ڮ���n���+����qEd���g$�4-(	�����	(H�l� C��[�.�bs�o3�nRw����]� ���w,�U�b�v ����u�$�%�H7�P�S�b�-T��?k�b#��8>�b+R,�=1�ܭ]�H#W�`�;p0KS��c,i&Lډۏ��ɩ�c�q/٥k����~�.�]ƞ�Z=v�w���]%�P�oh���B�}�t�ϩ�'��6.[��������B٧�)ǰ�F���9*�)-ld8/����^&qy�͂k�qt+�+o7����a9I��]i�Yy�������P�i�Gge~��ƴ�ut\���_�~���l�W��c�Uz<��/�5}��t�Ǿ:]GRw䶻����?Ho��L���_�&9z}��if�Z�t�����[~#=����^����G����ߒ���[Ճ>���������C�����z߃�Է�������X�����k���l�hOnL����/0!��a���q��i���GXۿ�\e��JY�7��w)�S���p_;���� �~�ć����vvX���q�a��A0��.2���M�+JP�<�铽mx��z"_�����DyF�2^�$��!Q �G���]}�* YD��,�"̲�<|IpLhh.�)�i�Z+��/��`t��	'� �z�n����O�L�l%4el��I�,���#��z��2�<�~��]䡇�/κ��_ �������~���!���ݼ���)'����{�`V����z����2qy�֝\���r�
㌅�,��0�g|���P���S�~C�il��e��b�L$����jɺ���dlÁ�66(.Lv���z�2ȩ�ڸn>M#�Ѽ۠g�5�����^o�B�J޴3��f*�t̮�o�ב����P��f_A�-Ey:����[g������ܔ�y�XT�?���NBj`"���Ri���8�ɐ�͟�$я}�0pH���'�M�`�S �F�Ř�{���#���������%����3l��o�{�F��镾ԷՓ�]a�����|]�8F%a�b�O�B���P�}�k���^̪ ���ͤ��a�_Ae3Ht���ur6R����լ�����^��|j�G� �Qt.?z�x[$��(��VYw�a�@I
WPp���muKQ��$�c�}  WpA���!#ĭ	�C�c&��"`Bl�uLJr?�`x׎��
���M����>�1t������P�v�\�6_O�_Q�Y�r�pyFwq;]�_�kR�ϯT�\:M<S7��*	y����#�����j���tun��޷���B2@4@�S�ui�� g|�{���lE�S���0@�h6YG��/ae���w�T<���U#� ]�&<G	C�7�3����_�y0$ӃHN��z&Xu�9t��Ϳ�;��-������ỏ��̯�=��)v�'�z�z�s��[�J��XP���Nh+��G���;_��a�s��t�r����j}cǀglp�+}�P_��'��о���#I�*�r�p�J��\���\4���B*Z���V�9������]	��%�iʻ�%���Og�ſ�F]	�_7��T~�IrRTn�c��{0��&�6���� I(��L:�nQ*���*F�2	�O��=J�����S���Ƥ3e@H=��7�l���� �����'P�����}F6F6�,��g�K��2��x5� t@@��_�&PJ�~7v󭑻��n�wHaT4� ����'ZEe�q��4�A&~?�k�m��,��Y��Z�?�����S��@�dV,�����4����n�(��+�!�i��M��^7���0����>M�D�S߀�i�)S)�w�5�E�"3A��t�����A$�U�ȼ�bJ>�gT��sc�۱��s���o��d�.�b(�O�����
���?A|��-J/��$�MHih �C0�L�%��VN��qT�d�X�Z�S�B��9@+X�j�_8!޴�:�?3	c3F/������68��I����v!�I����>�������p9�6:�+�1�i#֐Z���K��xh-���due��_,��" s�	���Tũ���Ծ�8�Fh/lW�+�*�U��OCn������G�����$��Ⱥ@Ȁ9�H�%;�w�hC�"���6��V�����0���7W����E�	f�r���7�jh� ��[����<�}�h2�ۢJf0� O| �Y��C�V!Y�ڑ=L�ڗ�aK����`}����~l[M#<Z�|�����_��WT�|�t5C����}��d˰��Wԗ��/xq�������+��%��e�ы��r���7>��0�*��s \��!U����6v�&F�"�d)D݁'4mQ�ܧ�_���w����w��F��l�<�u�S���D�x�oTq�Yk��tP?&V�1����N����5��t��1z�(��"@�mv�q5Ko:4y���P����:_��*��޵��Uze�,Hֺ����}��0X<�^������j��R��=Lt�QۘH�����pG�p��i�~~�_��ͻ��߅�����y�|��*_y++Ev����UIl��0� �J\��x,\h(��J���;R�ho�|�=h_Sa��g���	�� y���Fj�LWxG�ƍ(M�R+�tCyJ�hu7cH�b�� 2�I���hJ0�Q����~6�l�<�
�I�ȜB�a�: 2j͕(��b��c�Q���Tڿ[����)�]��KIS�ry� �y��O�?]�ob ���W5dH��W+�x��|���<�ٙ64�Z��F��nl?��H�[����q��?�)�^�ㅾ�M�� �fx� '���#p�
��Ƞ�J>�	s��$��"b��j�ۄ���P� U^Q����$���E9��iK�є��Ǉ��e�zC�n��O�SHP��ܞ�?i;k��^��`���@!�0���H��d�8@�#V�6��!W�6�m)�wKI�{�	;(�l"š����)�i .�hYJ�ɰ��>zG�D��!����.�?��A�R�]�e�e���!���\�ѝ����sãL�\�1��a��6����|Xɸ4}+x5��tg)o�ME�B�q�:�J��>���)������镺�Y�*J��"Ή�,�Hm�;跜��Ă��3Z�z(��c�!���p����h�v�[���N!3΁V�D����'t]u�jzI[llA][���6V�����l�q����̆V��A�BVvPvF� �����������1�N�if�3���܌b=��}�|A�o����o����������	��?]��vV}����r�5����ڸ|Mҙ���v�؝��J{I;�gY�w�L�mۆ�
�S5܈9�M
u�ߩF�;^�B_p2s<$�Z����
����D[�Ў�����9�_�U����wI�,����U�j���S*kY�ӞCc���r��8}��0�)ir�f��r\�gt�:3K8̋�����N���-Wk=K;�h�fk�p�T�R��4R6���+�K���:`�mX���H@�Ř^Z���c�mc{�1���'��0�Nښ��hD� H�=<��������.��;�,�wy�l�~��K��g;~���ʏ�� z�4ȕ�:=UXޕjQA8nz3��I&�u��`�i+�q[`S!��ō�	n�%ap�P"�/�����k!n���º�s�Vd*�$���i�AtC���2�2݊�|b���]18��[��3���o��C������#_�Ⱥ��	h��N,G�O�c�����D*�h)p�F�=��J�JW�F�Yx���/��P:b�KA�%-��~-�>q�Y~+�n����]����Q�Ԧ���M	�i�8B�.��Vj/�#�3������mb���@̽��k0�G;蹠����m��,
�d�@"����n�����΀{yF7��'z��m�ۮ���'���2$c��j�*xЌv9��$Я�P����� �׬�!���j�Eul*����<P't��|�G�m��j���i�E'������͖f���q�����@�Bi@l�x��@�$A����/+�E|~�D�b��9�X�1�g�jQ>����hg�vd����G)8p��E)�O�.'8�E��K\�0����%b�������FنHk#�M[��S����O�!��G�5xg������}�2�JA1c�
�I:U��9�0N����xg��Sidd�����'x$�{=��[;\g���̤�4��8 1��X�N%H �w�/M�(��wD���׭����k/�^�����R���Cj�}=H#yĺ����426�^�I�`�ꗾ�t���B�M��Si��S�>a%~ۋ(WO��::k�?R#e�N�閻���6��9����И�����m�C [�Zc�;��1��(�� k|ON�"?���GyF�!��8ٵߣ�2>D`��[y"�E�<��ihWD$�T�֏����mN�9� C���@���mT�iO���~���.��Q��c[S��b��%�:0�;;��!��$�۳0�#�ë����/���r���o�]����ߕ.\��ʹi�pz㠠��E<b<ņc�ػ���f��~6MV]�o��\J�v��W�<��x���-iK~�7^�so|�����d�[�K 5|���`�w3]���ir���Ȫc0-sE+Q�q� *]��Z�6/~��f�S"� 'A��ܔݸy���}	����:Ka�\�ك�*$��Θw$ ?-�����'�MM��58r����u�vm%>�n!��{ً5w�%��U�"$Jm.�{��`�u�C�~[�q)��AV��C��GbD���ͲJ� W,���Ǆ���H]�(I�~T05O��6�hxL�\p;�;��I��/h��f��~�ǖ���~,-{ɤ"�X�+:ET��J�'�:}��B����
��ؗ;����we�hi�n�b��#�HB(u!��k �+��wk�&'I�!P<IsU~�?��%�Գ�Q�#l4�&��G��n�ǚ�Y��a�P[�N�`ug[s��&�1��_�ʊ�t�;�у�\�OK^�c�{��cq"��\L<�􏀼D�ģ��9Tǣ�c�k�+0�ۜ�Q��X�dܤ�;��d�@'7�l$�Axd8��s�@��Z��N)T�  @ IDAT�+p�iկ���c�ٜP<Z�z�
�3�ї'J�3F�κ��+����L8��g2D�������*G�->��}HM��G1X4���!A8�1�c_����Z��'��U�%�MƔ���'''�יO�1}-S$�"s��6���*�C�A<��b����<'X�j7	�����7��`Ԑ1�W��k�^%Lo��`PңL�gۯq���� @Ὸųi�h�rq�Q����2GZd�	,=�	M��}ܷ��Êݦ����q�s���]��8�q+_�%4��^�d�P����0�!�WR����2f����Ng��_�l�3J����\G�:�ɇ�	��	Z�����!iA5�e��cWI��~.�(�d�ځ2Z���R?���V�)�f�E��r���������q7�4���:�_ezlGoo2��9=؋�N�����i�o��ih�ȡ �z_FcH��{h��c"P���Vb�r�t�18�X2Q﬇Ď�"DD�p�͘���Ejfn9¥�:�nA�X�$�g"(�Ae���[�����:Β7�;pW4`8e�`���Hkl�n�	�m=�Hߏ�9�q���D��6g�����癘���f��	�OL��	�3������Lgsuc�ci~���p�� ��lZ�|�~���`pn��BE�$�xg�9�120����NB3��(�@z�z�c�Z���V�P�����r���	�텇�{��Y\;�����ϳ]�{y���f��-PlQ��Q��Xߨ���W��{�3����4\m���Ʌ^|g�0k��!%� T9�z��y:���	��(]�M�Y�rG|�M�㙞d�� ��"��	!��3�2�d���G���&}'�.���1=��$�*�oV�U�o^���;Q�Ū�K"e���&��@�����c�"L��!(@.V[�:(�GL��x�j�1�^I[z 1 �j�0T�+�ܔ�U����		q2�#M��/� ���210�;E�
��7ao��b���U��>��S/k �<� �Zd���H5�x��0��>/�(�Ų|�%���߅�uQ���1brl��0�%(��N9�������U{/�,m��R��BObQv����;(o��и�#1������`�~��t��?MgO������K�� CX��ڿ�A��>{5]g/���k��d�ݳ���$�PՋ�\��껒�a��#�hD?� %&�7�&$Q0$�9��:D����1<.߀�(��z�����w(��~��dVi.�ˬOg�/�D!
!o��P���R�	�������	��G�&�ET�࿸
."�2 �x��gl��~��֖hu�XqZ��w�w<���,5��~���� 7���F�8>���d�����͞�֋W-<�F�C���Q��Ҩ���ez�X�qo�[AkKN����K�����w��⬮Τ���YG�TKK���J#�)T���֗�n�I�!��P��t1�D�yI�A�"��s;�no��^��R��Q=2N0��[o ٲO�-�
.Q$�7[E2� �9���@�$�F7�s����^Gu�;����Q�l[�;ظ`S��:\-@��	%pC)�$��	B~R%��lllc�^$[��tz������>�t�s����;�����g͚5k֬Y3�[�^��7����G0���i6�y��	��s��\G�"��Qĭ���5�8w���LsC���r	r�w��LɚL�e�#�DIS�y5Ag����:ü�Ew$�0�
���l���~�,���2r������Brg�
̢�E�4��Uq��-�E��]ɫ����Z��T~�s�|�c���/�:t����jU�?��"|̡c��真�'�ޗm[ۙu���N�c;�6�o��H{�5;��s(���񉚞�]���tv��w�5���z״a҂�ȣ��_��~��"c0��\�)[��-��i�C`Xkng���(ֻ��J˝AOj�^_��^yK#� �-������P��V9ۆv���0�}7B�{u�a�wϧ���<��!'����g�������pӕ߾�n�\i'#�c�p=�LJ�wy�3�HO���l���L�N����~���2�L
���X��[� [@쩳`��poP����C�5�M�"���J
�=�N�Y���0��Ƒ�Ճ8��s:yX��#�Q_i�+}��e�mjd3��
�E��7g[�{��e2�C����qMzź2�P�BB��_f$&�XHp���:<�ä���OM�B��)m�esJZ��ax�e� �s0L��N�_�E�L�J�-�6(Q�a�G*�T������g�ˇc΍i�#®�0tł�G_�)��Z���:bO���I���7h�4R)5�O�w�j���%m�0A������f�9�%L��̓{�
Ɇu�pc�f��P�"��O�������0�-H�6n�ȕ�ӱ�i��9=���BB8�DZ�i&�y;�:c��쭬�[��dg�܊^����[u�什9t��
�p��ʀ��kH��K��V��6�T�7}1.
f�*��d��"� VQ�ŖJau��"1����T�!r���L���0�Q%�u�0P�����XmZ��Q�I1�ˬ1>��:0G���:1V��T�nۚ>-�	��1$=�X|^¢�'��WQ�#�i�[���rϬܠ�3�J�)�SV̼<٪���p���Hރ��vj8��jvS�f�oE��>|�iǎ!�O�������瞋�0�eBj\N�(��׵q��Ӟ��t�Y= %�a 8݅��4&��De�, ���!����v� '� �ϓ\S"Sc�K'E�� �z�X��Q�f�f��3��la�U��w5��hE�@s�+�D��_�rs�<�$Lrheَ��+�OOy���6�쌤���e�.(�ՠ&Q��ۿ:�U/�.�|��7� ��PD���/�`T�]Hb��A�D	�#���fP�Di,m[d2�/g͏�!`�O�Ic!�G�x��o_pE����_���{u�"����	��eX���7e�u,�Y%�e;�:�,�-+d n~y؋~a��������g/x���_����I�M�|mO�J�3������j�c��7�9=�������=���y���lڿ��骫�Ho|������W���i��O~��i`����G��\��;��tW���:���0�4ao*�I}�W�\�*�3LZn1q %~��N�3L��i,^�O���WɃǯ�U���,����/yq�F,�P����R/�[|���!��`u��sA���q���#�x�ƫv0��N���g�e:�% �m����1�E(]�Z�T\�o�)"B��'+�!�|�E>C�������'�bXD7qGNЧ�������P(�����)KF��d:F����l<Y�E�HcY�Z�9���8�j��@��{8-ƥ\Vz:I�~؁��"i�k�����^� O�4.��W�.h�(X�G�9	3x�@�f��f��>���a-`E;X�p4Y��Ƌ�QG��g�D�^�gݥ'����G��@�Y��PR0;�
��2�#ȇ����m��7�9ByZ�1D�v�{ESj�!+��3p�r��l!<L�K��(�	��F�W%[���3Lb��nxG�����1��||�U������(/v'����DN�;U�!Q>q��b�#A��`�*�oK*.�m��|�/�T~��(�r�x�qY���^D�ǫK��mM�)�� �1D���k�m��Hxa��fg�rB�q���^�:�ʹ��fa�m�����m{��ì^��f��k}�wϞ�c�6�]B���ޔ�q���y;&���?��'0�3��Ps����5l�=���XLpz��5�ۻ:�6�}-�I�fB6�x� �" ��!�
��=� p$�D|�i��E�[���%^O�4��N��,\�J��O�zd�tߊ���p��j��M��������M���� ����̢�RǢ���=?r����,˚�l7/q�����X[���֜����X�U�CzD0.?2S����[8X��3*�4Y<�Br(��dw7�f��n_�^��(4���@���d�^����0�����O>��W��Ǖo�+���e�P��7��ʈe���gV���+��bX��ݺYO�. #"߼�e8�D!����Z��JڈZݟ��������ײ.�["	Q��8m�M���*���엿�e:��%�`,>����O�Yz�[ޙϷ.f�����n>߈��SH<��zۆ�|׆F�e��І�ap�N��G��|B��?}-���xh�]��\i�Jr�l�} <�Ѷ Hu 0�;�i���8���ʸe�<�?/��0B���{��/��>]u���Դ0 ;���U&���-�,�Ն��o�#�^�\p�<U�ȟ�8@o��+�0�E|�scbœ^���EH�,!V�'#��	�'1�y��@�t%�#���`i��)+�_�!/�� ��|W�ft'��.�3��F#8+�}�H@yv�!zLFdT��+�ZO1�l����C�|�;fmt2����c���.�*qP��+�1
_�(�i����c&
�9p��Y��`��B�o�"��%Y���̓9#����0q2֓?U	�z��ݙ�Q[�vт�aK>�W�|k�zIp�n�b�"[���h�zY8������7��&0�llf!�]��D�����,V�v��JVQ�F������Q'�B^R�i*�O�PP�0��������,*��;�ȫ��O�/ QdTyf�4	��ޔ���X��V2rz��o�I�L9�X
5s�t<����Y������A�Pypn�rr��C~�5�������o���ZB�Cq�9����,�2����/���l]i?���3��.�q~�oZ�;�����A�r�ݓY�ԣ�RJO�xG�o�+
��NG׉�.O~|4o�r�8 =,�ql��\P�b��C���.f�x!21�o2Qig �"�e;+�X�x����ci�葼�k=}�$6�Xl�ZJ�䐜�dK0(�i7F���d\S��2.���`�%�$��l-N��{N������㧤��{ �o�6m®Rkz`���x���U�(R9NO�fJ�en%t�]˪$�ޣ^XN�㨥=.b�������|b����ij�)g?��p�� ��7oN�3j+a[b_t �����xYbU��ڟȫ�,:��J�ʋY��4��#��cҮ���Υ��A��\|쫀�����83�Av <�
�rz�c.�E���_���엷ߓ������y�����קW��Uir�`ּ�4�5���ǝ�.~����wܡT�X�")b<t|8��G9��c�p~�3���h��ً��\z�c�T���=!a��߯�-e���j�B�r>�9��&h��0��g �I6[���G�2�|�`q�dV����t����*�ʧaU�갺I��}�����/�$��^�^�9Y܅�r%�R��!p �6wv\�HA����~
����Sl�]{B�ղ�2t�Rb;ϤALH,�\��p �g�a�@1�U	6>�<�*1Z�*G�+�N28jŮ���(L�hn�F%-�o�$�~�n|�H*#"����3�	����Em*�Y�#��Ș|A��<W&��<�X�N���8̉D��d:.�vp���������t +�\���V�f�踕i�~�>0�jr�kZZ!\�����I&��b��c/�*MR���c��P��ţ|�FF�-+'=��B`=}C;��ÿ�_�x��❣!��~A[�����@��2:J�P�Ȧ�-rM�pmw�,��a=��)[I�<�M�b
;,�)�	x�̹$jhF5�y����!`]��O1y��6.ha��Ӽx����č�7õOS��ѩ�
��s4��ǌ�"A�2�ѣ,�y!�T���\�I�\!@u�R�����h?�1�[��-��1�PL��5ܧ2���`V꼲�"L4��A<o r�Q�x���'E0H��N�F�S�� ���떧S�#j���ƨ���ݸ���u��l۶M���,R����%K��yR-o�t<�����á1I���9��[�lm�iA�'?�~~��4߼�mA�k���R Ϩ��d�����%��8@	��#^IAU �~Ev�����<3?[Ӂ�[�cG�1�xk�U���`%���)Pِ��(Dwd��S��<�DO�5k��@ y�ʠ��2�籒ٛݼo"�����a�e�FN��-/���ǽI �{��$K˝w�aL'����H�c;�UDD�;
�T�)d�@'8[�{K(}C$:z���؄m��b��I�$ Lf_�U��t�E`����P�E�����d	����_)?b��U�E�Ju�z����H�J���M�?�Dq�-��/�v�Ռ�G�����ݜ����Qpg��<5�n����/���رc��ml�Q��	����E/|F���|SuT&8���h`�Їe|�����ӧ�����j61�K�3�;w/o����l�؝_q�%ٷn�]�`�^�^C��#=T�n۰5Y�����M'}�'?�(����)��,��j��2�ߍ��[?]u>��Y����g�b�z5�Y'�Ǉ�O|�����zf������ŉ����S��<G9]&�k�o\.�{HT"� �+�L{��[�?x��hx��}�19��bƭϬJ���'�F��!��n���4�L��$\��a~�u�T�ʅ�R�j"R�p�bE.*�R^L2�GW����d��T�5rW*;EJ8�=���A��2e���(��p�Z	��l��{&ȣA&�D;C��wt4��#c�ixdiEM����{z���}CwA%q��"t��[�%��[�λ�b5��1`=�1Q�9!#�q?��ٽ�^u�8)�驟l��=�V�Ǽ9��lW�5��vڝ�?��Ca�����ȾW�R��qI���'�LϢ=to�:���y�j��1(N��U��݂�ho�PhM�lK`�%�7��~�E�u���������	t�Z`�d%��n�q�D2�	&�SM�s��:N�u�@�*��F�Ї�E3�IFm��"�<����w�V���	��e��M-]3�Qb�1QTCz@n��U����\�7�ء�#�'H��H:O�yQ)G�����d���\�rح�)h�-�����6q��4qb�v�%'0��k/FK����ผ�.�S_��c�up�����.-֘��%�8=�+U@v���	<�յ���1���#�;X<8��EoWo�=-p���8Aȩ��ǆ�(س,޴~�x#����9�ޜ�{o���k_��ǟ�8p(uq��i��ÜSq�R����t��U��~{�y��P Vay
.�����4P(E���ԟ�7���9�;�`����7������o/�n>q��el�]�	
=��[} N��G�����,��yŁ�e@���@�;8"��v�jv.l�?JW268��y��u���sDjD��>�k:��/x�S�M��5cH�f�����˱y�Aٶl�`�&U𭫖Ke-�2qZ�.o�}V%-Ɠ��t������+��v��hw�3�n`�A"�<\`�,x(�����^����|�, ��dK��Y��X�U�E�+~���N�����e8��?�I����K�:�e�A���]�4�A	 H�`!ń�VV'�5��斐L3O����Y'�ן�=N�.�$a�������4�~}(u/�;�}���'>���5�zq���>�o�r����A��%��gW��Ͽ�H��o ��yV��md!063Vs`x:�o��F�9��r�ƄU{4uS��lb, ����-���6�G�����k�2]��:��W>W���+�N[�W�/�E����2/��-�O�
�� `�\1\�u��Q]O3\>����9@$S ��#�b�7F!_#Oh��y(�(1��Š��Z�Jᴾ��Ap���� �}V*V�)G�By99��\yG���K��X�)~�,��K���Q��o��tJmV�ު�42qAEԜ�[L���b�dV��Ī�f- ��Ht�jev���N�]����%�H���̧Q�q�&5 ��D�:����O3���s	@pP���Iʥ�ؾq.5SL"��zQ�8�Ƅ^K�細�	@�sL�!Cp��ہ���^Z��i�g������& ��$��0�Hu���f0k����釥4�����,Q����J��j���	8BL��`bݙ|c�*(6"R�N41���H�6ȑQ�rꆸ<��x��+�n:0���}+�9������j@t3K�����̑e����D@b%/���$�3�`nDװ!�r�NR��G�Y9���ˋO�'  �,����h'��1Nb ��8e(L8�J��%�2RdĜJL���(�	���~�v]t��$і�9&=��|Z��.�s�r9B���q;�D��{�����<1{ L����i����ȶ%�""7��01��O��y\H1=���s9�y|��x��g��sБ	���1,+�Y�6x����ԋaH�@ �c��3a��O?Q?����>�8[A�0�s7���S�м&}������z���s[��ؖ= ]��Gw 1��Ssp����ǳ�3ql���jys1��j���u�c�.�,d

C���NaA�����ZM��+	Y��o�"*a+�����O�{���+����v�, �f��ɀ%���D�u�����t Gr�j �w��]2.j�H��1)�t�I4�+99*�5 D=��:@�%�J2m�[/�x!+S�;�c]K�~d�X8�#'��zX���6w�[8a��ka�P�W�*���UN��*F��{D�W�P���F������~*�x�gu����q#o��i�����Ө��b}���`���N�	���VLa�l��i�)���{�K��.ۙ����A	s
Eʟ�������s(�aj���Z�i`�����7�V:x�����1UȜbY�o?m{�u�2@c1�p`ƭ���{8�莻EA��g�r/w�o'�+���8��i��5M���HY��0�>��E;�_V����w�KW�W�U�Q�Y��YF�^>˸�S]YN�u��7~���'+���L!�@!:�Z�9�A� �nK����`�ihA�,�`�����D!�;��9�%֫0Q�~���2�G�
���E
�W�v��1l��K�x:�9#⛁�4����E�+��x��cj�z�-!E��	�Isf�=s��uf���IbiiEk[6o���+���՛jm���>�'ld��g�s���<JB�  sSX?�T���LֳnK��]=m��p�6ʉD���F�&��ST�oH\qj�EEWH$�hL��PxF,�.A e��Z]^�~�t�cn�e�}��3\��5��s�?��9ǔBR5��R�jӤ��`��w@�!L�\��LS=�w��p�l��GX	: �k�$� ���@�U���KD�2U���Chf���^� ��mu�s��JlzL��}S�ع&�&����
|):���w�u�NȐ��G2��`ʪXR���U�B�;�_P��h��5���	&a�n�����U��U�+9�破$&���[J C�DT��*�e��9�5�EhW�r�&��3ud�`I��:2ExML�/�c���Yb'cj��3^�)UA�^5"y�m�D�[���?���,]����$�y�_�	a���Jt�&��R�$�k���cHk�2��D/�������]e*����L����t�*����Ӿ�ZS��0 �<(7���(��`f����z:6�K!��p��!B��w�T�5�"܃��X#fL����1�fP"CA��܌�R@5ΰ�)+��Dq�1^��<�	�tp�hrl<��`l7�AY���et$�iC!H�\1�T��h�N��
V�ZM�b���'!�S�洃j��"�ē1�g0�J��迋!pP���E �6�m �Z*aκ[=�G��M&O����6!�
R2c¡6��W��[�E��5��)���|A��С&$'*��g%��b��t�]k\Hl����Q��w�-��� �8e��3��:hY�+�C��cJd���:�3�#s���,o����:��;�,��/�tڎ�Ӯ];f�R[C��S�ݑ�<��w��_R��xt��=�$63���>#�b���w�1�Y�fS��9qڎm��>��{q��T�[����!� �8���d�m���M,������~�0{� d�i_	����W��_�HDRPhU^e�j���W��y�N[�+�e��8�����h쾇�K�`8\=CQ �-�	䙼\qu��ӈX�y&P�+RQ8�z8`\ACK�&]	sg�X�Vd��`��E�~RTA�"/�^1�� �j3�F�ND�4�1#1�)]T�D͊�7����RJ��9ᑎa;�O�������Ǩ�4�Ǜ��0iʆ����4�*�����G��gc`8�����5M�d�mD2Bb�8�rs���2%t�Xes1)�M\_Y��f �۵!|�e�~̵��x�$	�+����Se1a�D�#�T@% T�`zXI৤	xA�Ѕ�����Slm��+K�䪥C�S���5�e���y���v����aU+R{�S:2��D�Y5d��9g#k��@&t���c��p��?#g��?�&�l،��R0����]�L9������9���j<�ͅ�R�%0j����AKl�r� �%|R���'{����e&�i�	�a��`Ҹ�H�ul
�������U�A<��5Ԋ��XV�8��6gy�M�c0���ĘR@�Rj��S�~ �2C ���U��8��y1��m�L3�C��8��$y1\�F]8t�=0&h���`d���%�N��XP�Z��!U`C��&P4��{�zl��⡵�IE=�g˅���9�7C���h��ET�t���(�hF\� ���_�:���t$�k�#1�AP�3Q%�n�	��y����GIxYw�uQ��-�G�+RV _�c�����{�"�!W�a�N�"���2�%E9�]�@��������u-:�r�|��Ju�G?�jE��U��U����"N�j��ٸ��Q*m��"8`%�p���-/��i��qu���s���I��S���8�T�U����e��=d��z�4EQ��ZJ���bn�μW;��wYf4ni��? cZi���3'�ҿ{ɾ��_��z�mk�ғ}& �`<��k�΍�K��t��}�;>���_����%??�ز#��n3�,�1�1����4t�����g0�`�����Վb;���39zF!i�Xe�������2��K�ӛm8@ƶ)\�{�#����[>����`qK?��)Ӕ���J߫ê��v�i���u����zѱ`0�c��c�?��GâL�DtJ��1����ə�*QҸ���*#[���\�ǊF8[vQ"�b����'����E\�]%� )� L7��Y֘Ej��W@9.հxu�ؽ�{����Q�4=>B.5�3ԫ�_N���̌�T�˦aВV�=3��V���6`��-����	��L�nG�n�q����yl�@��)��H\&󥬽�l]�8#层E�!�1�G����ʲ�v���:��V���j��SH�S�^G�nA�g���87���+�f3޴�J�%E���mg�\�@K��n'O�-�R E"%S�FН��џ���5{���S�^�8*t%��>u�IRZ%��~�+_���ۛ���w�zt����Mi|�R�bR�@�aX�|�������]��N�abċ��
bR��ײ5���<��*p;7F�0~	�ż1�:њ��3�3��(�7!�j���⹖k�aR >���N1��G��~`��s��m��m����mB�M"�O!�r����tI\��	R c�:��s��) �B$!f��SN��*�$���9)hH8�`ظ0�ѯ�!����*+D2m��`���i]�X���=M-�H��\q��̈JƷ�җ��w1��$`�)�x���6N�4��+�$K'Y`����ҝ>�#�K	�����J	"*eƸJy�N��d���R�x���aR�3 ��(
l���t�ې�
o1�IJl���=�?2?ʏ��P4��3�ҧ��WQ	R@'��c�qD�ȃ�E��"|�s�1䉐J�F1P(!ɢ��"�D�H��5{�*V���m(<��`Db���\
���EZۊ[I�]�G��'
��K��F1�y�_�]�/�։��|�
3����MU�HFܬ��9c!�0δ#6â�|�����t�w�I����[��>������K�8��G��|��	��mJ�X����(��g>�o���Ƈ��Zl�-17�rZ��]��s_�G��u���Ԍ �?�r`Q�Y�s���^;I*	������Y dS�U@��x�����ӿڑ��r�﫿��_u�2�����a>�+�T?��,�˸��5�� �>�'�
��(��e8����؄��@Z�����h0�t1Zu(CdQdV�dCPp���A�hE�4|�P�sŁ���KJ�2�l��?K2g����S��-�	9�j�V���	NHa+�s�ػE	��X��S*�vW>qK��id�V}�vT��𑐤�p:f��sۦ��ȑc������42:�Ԇ	����	l3�u6v*]r�Ks��ٝ�ݜ��r}�:����c[�����X@qT��2Z�mikOx��h��K�`���!�X�����U�& �Q�1?�U!�q+�?4 �e,�+ήG�����ؚQ�mjkJ��E�G�-�����՝�0�(��a���&�M�0�'!�`��Ǆ�~�ck�w�I}x�~�"g�ˬ,Qe<��b'!���ck��K��.K7�zK����S�**��(�S~��3��1
�)	a����B�����+��C�Y��� V���YY&��!vvz��/X&�˿�&w6v����!t�&��?���%���q��U�u��b~�h1#�A)�|�',��b~�)��̟:1�Ջ(h"�a.�g�q��w�D�*w��"8�t�yQu�Z�W�:���lAe�4��@�\��i5�cPV�7{���J��D��$�1j@��F�<��e���<y3�"�!:&|���V����^��+~�T���x�K_r�J|�FQcs�}�.࣏yXГ �E� %�_�X��-�2�qH%>���i��4�"F�E<������)��b�x�BY�2��dɘ1 ܹ��6�.OBC\Lk�E�[�)j�{�?jC��-�l��pE��H���O�;2�o�F[/�
�.�m��Nz� �=�I��Z�W��a���ǚDj#�f<W��̗��q�T*X����/\�W|��_D��	�W��d���V=��Aϸ� �^��o����O�.xF�8ɚ���,T�8`��B���-q�UW7W˰�}�%��l����ȝl�\��m�h@��{���R��}ߟd��R{7[��?�bo|j:?x�b!O,8����уن��� �
;6oN[6�Kh�1��>� p�iIX.�{2�=s�����+�l���g��6��]V���`���2^�G�,�2��Ҕ�����N[����Ϋc�����]���h#��񅌀�- ��%vŠ�fa�� �R��bhÙʀ	p���F�A�%3����X��J�;��^����y��O��&}����8XV%�+V�������ْ݇!!��r���hB�볶Ύ��Y$,f�ɀ�?rK/K\����D-!;4�q��0v� M���^�����SG��.DX�Ś)���CGS�X���QVCV�)>��U|ie�M!��T��V� ���!�6�l� s0��E;��8���N1�&�~!kF��mki�� v�`x��|o���`��&įާ�z�mλ��qd��l	6@�G�M��a�����C�Zџ��W�3��Q��*���7Fft� ��w2r��l��XB�pb�"�i���(nK7�|zHcycK[6��}rl,[b�RH��R
9�w�@�33=�}�|r4k��h8����q�N�s���ه�J��	/�T���2W��PTqB�6��U���ڱ��d6���[��F���ҋ"/������E�h �sxs(1Pc�z�.��?7��З-�M��N<��5c�o��d�Ȇ+S��%+|ɕ9^(�_!�`�6^��8��*j�niՍ0%?�X�������
�J�0���<����
s�*� ��q�9�s���Y<c���SVƮԋ�� �j�$F����4%�W��Udf�Sg���Uޣ=xK(����OO/������QqrA aɃ�XXm�-22�x5���J&ENe~�SV2ދ6i��S�'4۸t�Y�~b�*NozH@'����֘�;ǘ���m�آ
�)� �`|k43�ؾ�h	��H��Z�RJe�~S�4���idx*��	�h)��DZjQ�bAJ�Q����,θ1D��v{3`J���o�?6*V^��uuX#UoG PGFR�h{�����&EV�u*���(kUX�U���q��*�xZ�J�H[���gx�*�jp9��=9�<��C�Rc͆���%����ϯ�Eڱ}{��w�5mX��%���b}v��L���	ՏE�����3���u7�NO~�vnf@Q�*,r�B7R�V��cqV���w�}Й��<u������yw'HiϾ�C+�[�|e�N�����}�dW����Q��䀹m;ɿ�^����W����_�fu���y�[�]�+�N[�����B{#���)"��G��&Dŋ?0�8L��*��Xq�(c���Q��ӱ�� wZ�� ��H�u���X6=�Z�M�@1�t4"p�4�� .�3MC��j�W����ыQ��Q��$6����gmIglX���n���5H���ή��v۽{���֒6m\��h�� ��{l�|�����n&����c�g����_K�n]��8����g�k'�0
��Ԓ�9z���y�#���V��Ng���tvw�:X��'	a:�Θ��I����o���F]�Z�%�r/�S*�xZFZBK���v�ï��\��MQz�z+R���|	cnG�%��/�N߹-��*��w��~������Һ�~���4�tdӺ�4ttOV?7�^�ҫ�$�=|��;_
`GrV�Pl1�Wѱt0w��' �ѕAX���7��0趤�����9VPw�ɾ�ѣT��m�Հ�"6�G�'X46*���!�C'iv<_�۞�ߝ7/�eo�o�����_��o��`V�	�2��NPr�Wؖ��)J���[�����L�mg� �G Z?��@���~9Ma󥾁a����X"Pbb�bj�6�rP�d3:q���F�][֦��o"AL�'��[��_�%ǘ@O{��
2�� HkI�Do������ac�ԙ�3X���,-��̦1���-���m%	ؤ�u財47zd��ʤO�+�b^�������*`��b�0�<�W�/,�Й.��{1�F��^E\�)Z�H��T���۶�h�RkH�et"� O�P�q��Y�W�/B��c�T��j��U����>��O�W>m_�~�ꞥlu��M���ɊP��EA[���[��i�}er�2�me卼�"E����Y��{"QcVhk�Y�O_>�aÕ�C�ھ�ԚL
8�gT2��iĐ	8X!�J 0��/�$�.<�%���!�$M�R8M�H`iDf_�,�#>�������E��?��*wr\���J}N�T�;�S��(����a��.Nצ��×��w�<mH�����t����H��������}v�R�)�FG)�CCS�sMM�v��?�ɬ���i�i�i`[j���M�q�q��7e�����C�9Y_�B�mń
���oݒ���N��������]���52t�x���O	�h*�g�l�I~�wu�~���<V?����������y��Sf���e��O�֩���&���* �r����am@�"�[��)�_+�.e�yst��:<�N%�t‪�0�jƆ4-�Yˡz�'�)�����Hd	"�����  @ IDAT�xu<9��k#qQs|���H�?\�A!ոk�����i�/��7?5�_sV/oN���0rAV���y���X	���.��'e�����rk����s�?ܝ�Z��F[gv����]�~��O�Γ@.c�D�*�i��(iym�-�Vy3�k�2��w=5�񎋲o������ݒ��mLM]k���a�Eh��E%���/q�"���ɱ�é�S������'=-�~��2u�V
� !@޿XL=��d_��9�o?�/i�+]]k���,���|ij8�ȇ� ���-gG2��uw�Q���n%V4(?ѧ���r�olF0v�����´F���N����7�7����)C�|br,�d�O�L�4t�r�/g�#1�G~!��P�@�S�O�"s�gv�v,�f����/�Lk�j��N���o*bAw�1l��M^Y/��v����$UD�QT�F�S'�a��>uC�D��	Z��"�jY��7�v�헁�g���z����������v�A���;�Ր�瞦��OO?���O���q�%v�d�I4�VIS�{��H�w��7�qR�8�6.l�������Ԏ/2[D�LvL�u^d9��5صl�,��f��Y�OOO��\,l�F�(Kf�Ɣi��G]lyY1+E�:b� K쬂��LҶ�^���8&�?HPy�ҫtv>·y�L��*�.`&�N����Ԇ�X��ɤJ2C�P���,��D� ��I��G͊�J�Ň�(pw��o�F?ձͿ�P�� G&�(�H�z"PZIǋ<���zPo�׶�¬_%WC"�%p)��XSGG���ɫ�O�h�eD��8��f��uQ�S<t\�8VITQ;�B6RP��*��:&�!- �*�]� t?��l+�B�qN�D,c���ʣ,k�C��|�O?��m�J��[��|���'���r�UB�������z˝����fs�����g�|݋���&m��oE�R�=0������N�Pʿ���e/{�%I�O��M({�@���7M�7�������i�.vB��o�5=��P�s}o���C}��=�1h��Ѵ�O_�Ϛ����T۾�Q��0�;��bZ!U���v�o���r��O�W���>)A壌_�׻�+���}�iV����̯�Y�]]>�S�V�vE`
D��ݢ��)�5i �{�yGȗs���e~
ìy>P�Yi΀��++8�kj���;�L�$`}��%dt2d�Izpr�kcPG�����;�V�Z>�+�p�$��z�,�Z볉ㇲ~����~9�-sJ���fpA%�kn�E:64�=p�w}Mg�C�ї\�6�g\������e�Lg�A-�M�_\sk���+=�	W��.<�iq1�2�`$�ǆ��o�5?笳S����,�4qg���d�����h+��i�i;Ӛk�&�Kw>�?�r�Ӳ����ALO�˚�M��^��8�,Ͼ�ӓI	��x7���Lvڶ��{�vA���Z53(>�r�P�N�şrŮt6R�׽����{�vZN��]���������`�Rv�o۶�4���$����n�	=��C�O*M����#�T�Y�B��O�C�	Cֺ�
�M�y�P���lgrn?�׮Kp�@�O��6��oiN{G+w����G��n�{`��c�ܶ��mDl��D�^�ײF=T����V��n7/a���Uқ�����7�Fv�c��n�����mʰ� ��>��`�4�B�
�J�u�M�L�b/ef�$��f���Ѵ��!�S�p��@��8�-261�	�"x���P�d���'(�����G�Oi5�'_d�����+d[�_P{'��C��y֚lۮ�_+��S5�K�"����r�
�i�n�Gxe�����|JU%W^�h<ƏO?����������N�$��2�ʳ�4�\�2R��(�x��3K�!���"ZA9��y��'r��t���8�����"$����F?��q�I�4`N�9��p��VP6)�����5���_a&S��1�� /�E$���f /b?�1�vP����ܣјJ��wj��9������s�9���J�E���}�aKc1LB�i(suH�'Q���%�x�����.�h�p����	/2?�4i�	D�+��v��u�_P�����&&g�� ��ԑ���>4xo���ezꕗs�,���W��t��wdc,Z�l݉��P����8���ɖZCjcAξ��}���о���{_j��˶]g���~�s��se���Ѭ���{?��w���g_��N�v���5��֖�	��tUY�F��\���uڐ�8�A��]��I�2��S~�w�e��]��/��4���q��e���_�Wu��"�"=�`1v��$\�A�^�A8T���ټ	�@�7N-q����������}�M��M�\�<�}��:N��M���Z;U�x�|]��ņ���h*/��Ro#��G�����5��C�Z��h�sn3� g��~_�>I�f.�l����q����OK��p�f8��t�ӫ����KzO��,:� �}��}�S��R��t�LN�f��9�����đ��,$�nߐO1�\{��t�m{�G���i�s������g_�=����/��P�^���o��������{��JL���h��7�N��d]붦�YV��Wg�z�K�sM��.�K�_���7�����.�w�����p)e��� N��UG�
!�MQ�B���h֏kqdo�kC]����3ӄT���З�I��ߤg?����ũ>���,��^�^�������{��0�'��j�����L���6�g���6(��GÊ�S^����j�Um$Kl'�.!;�d��⸍�ݔ�6;;;cs���'����� 8J����vW5�c/�H������J�BU����bC��R���5;}MCz��z�[d	�<ȶa����ꄘl@?�&���gGJkнZĺ����߭�z��6�mk�cG������/9��j���\����8�fH��m��v�֧&���||f,km�/2NI��q��e�\@�Ĩ�����:X\�*�w�S
�����6�<6u�3�/X�N��Ǘg��9��E�KHu0��O�͉B8�H3rX�\�ܖ�7w`�S����)u�ćcc���R戔Ny[Ww6;=�}����:9�/=0va6`_!��k8 Á�6���fc^��ť�H�8����D����#
�ʨ֓Y4��r���'9�sމ`�p�>�q(�]8��ĳd82�@%G:����/r��
�4,�a ]��bIi{����D�yS�/E������4�c[
<��8OiZ���xr���-�#��8B�j��<�셓��1��c��6 �z����pE���=P�`3�FzVLN�l�F�H?F�l��#LRČz��ú�Kq�8�2)�*�(��`�Kc��T����x���;H���eI�!�K�>T�]}B�Nы�Iti>%��x��a�K�9�p!E�~2�N~Ojg�fgM���W�����h���-��|���_�E�����
����Lum����4��6g-[�������~0��/Ag�CEp�--k���N$GK�=m5{���Ip5@e����s�ܴ-��h���l���?_^�%����w��inh�ӳ]i� =�|zZ>cW:�1��F�����v�p�'aw][��g&є��r��ݶ?�p����_�w�%�}�W��o���J�2�̧�.�+�����Y�:�,��|�&��h�H;7l�@�#��q�J�cH�QҜ�ր�6]�͎�޳�������\���n�82��c���i�X��Ĝ�`����mw<�����m:46}�����&f�v���zDx-!r�s�T�a fg�+m��y�S��x��'{�|=��!ñ�ÓR��|��� �#H�0qX?}�y���t,��{��w��*)U �$�������?�>]�k/d�זi���������_�G��钳���`|n!g�φ��(`C�}^��6q�'�Q�Y�v�?��Gҩ=�K�~W���Sz�N=<���)�葰�b��28EbH"�Y�
a�<S�A=�&�Nn�>r�D�q�9���l%4���_��������}���OÇ����<��N��~6�y�� a��J&���ZiN-�L�\�	AC9]�fY?�npD�17��XUnn�&F'RM+����蜄�9+j�kP�w�q���ҏR��X��QJ;%�ė���;Dvݫ9$=o~����c�i����/ya���9u�X�b����p�_��-���=�Y�fb<�%ovp'V�㡽�fCG�u}�5	�-�S4=��uf
�SSܣ��Ύ�l�t �4�ӑ�w�=�k��T+G�~8߶�?{ʕ��t�ɚ�����L�p��6����c�X������<������0P��Ա$l���k:f�F͉.]���Կvs6>M �b���R���Ʊ�!�7�4G����H�<c7�vh��-0��ib��&�mc��<r ���U�K�эM�F3�׷�&V�Mm�K`J#���8�g�*�s|qՍ���,Na���1����V��S7^lY� Q�sx'��a>W�I\�ነJ�@� |�K��*=4Ml3��[���^����s�W���(!�%�/f��և��S��y��o�RtD-�`l�շ	��"��J�g��?�W0ƭ�b��E�0;�' *��h�T��4�w����u<=��eY�|Ih�(_8R�(_<1c�߼��U��%���%�1ߚ���I<c�E�E��_�2ۈQa��:U�q�I/
%�
�̸�&�<��%E�5��C���)Y�p*W⯧�����a���YFY���N��95�Or�z,��\ML��@i@���ݓ�T�
*h��Z�Բ�����Ҿr����ZrZ-Qu!1jL���6�r�hRm�{��X�j�,���i��n;$> _:�_�c���q��uXU�/�χJ��W�u5�`DHN�h''���Ps��6o@*�ym����={ �O�������G\|���r��ŋ�J����>p������k�=v�ͷ���Ç����>��{� +�o�֮�2�;O��	O���^rNe/��E���=X8VQ�<&*�}-
���1��sds��S��|��+����OI_�����~xu�x�%X8-t��]��KWWc�ַ�1[�+��p�hGڴ���g?#�}��/>���̿x�7ѧ��֬}�Io''�P�EO~+�I�D��M��Z�{���#�\@Xs)L��9�����K��8�3U�ɻ���� ���lq��&91��F�z[Go�k�χ�ܖu3H^��'f�`:sq����M_�ַ�u���fj�Ӗ���#�{��2A./oݺ��_�~Z�a#��z�-{1 mc��1g���ɵ��u-�g@�o��ʴ8�`�Q�`�A#�ؒ�9�co�eV���IuP��|�Z.��-��B�(_|�sd�	��֨�ej`P+{J\:�әoټ1�OYi�6&��7^zN��5?�n;�/��zVj�Fȡ��`X��ssjZ�\~��2?.��=��yoWK���鴶cg�y &���6���nɏN�g\�sk��gm���g>>�ڹ����Xl_{��食�|6>� za=y_:�/{�c/����'���)-ʮ���tƮs�������~���IQ�ҧ_�^��Gf��%cu���/?������9/x>�T:2<�����]s�-� z7�̛��?�0�ڱ���?I�7��Oy���W]���'�����g>�����d�\rz_��[��֚�v�S���n;�կ�O|��w��;ӹgo��nN�\���ܐ}�����7��]]�ZC�e/�(�r��Vs#�טĖ�$��g"a��7vO1'��y�"��8b���.��7��8�3n�Q8���.�'�ꭌg��9P��9�ܱ.f�(����xC�H�T�ȟL�9k_��(i}�I� O]l=�6_���.��Bb�{�Gv%5��d_�,������B�!�0��e�_ȣ̫�#q��7�,�AQ��J�VZ5/�d]q�VI��oʨTVZ6�2e"��,��TZd�Q �"�RipY?b�~V�æ�/��>�4+.�Y��Ze%��[iTF�����(�������tm���T�w�O3�`�������\d'��-���d�	��]>r)��-. _��r�`!�"�	I,$V&����D�<�8\J�iۖ�9E�0��m-������@�#��6�a𧭿=�e���ZK[6���8���`gi&�0��ۃ�&4|�!������ �&���t;@l�m�C�2���q}7�ڿ*��+���U�����{Ltt4�IQ��VX����`��nY�n�y`�m������~��߹~�֝Y��{W6�RiHz��<?���wܺ{�y�������59�x�b�9.�$!�@��@C�@����z$���A. Y~�,;��Z�?��۹��/"�`�����\��ZQ�9�@���_�^HJ�}v��љ8:���}��6qM7ľ�#.<3}�o>����m�/����M�� ���-g��e�=�g��Ԝ�g+	qw�3{���\��#
�1찛�c�pr|��Sd\A���ڛ�:��g;��m5�k�W����^N��8!� ,��4tq��8�����g��\���t����w�4�>N����Q�싯٘y�GQ[Pκ���G޿nsv����?�.�am\�֌܈r��Do0&��GyuXr�&��Y���)�f�!��f{��ˠ��aT�����i�f��ʪ`�J(o�:�8� �E~�
�!�Vi�n�Em0��5lT5dk�[�z\��!!z��V~#����)�F�^RoO���0tz0}�C�y��5��*-��7��?|S\���%�M��8||.�u	������ң�?;��e�H��@��.���pV���?ɯ�����w(T�`����0)A���r0C���bĠ�]��Ӗ��η��~ӻ�˜O�ԥi�|ء˹�2CZ�>����|]MS�!4�֚.��;i����=��e��/��5�zaJo������쒇��m_ǝ_�3����Bׇo����\�[͟�ηk���ʒnŶ8ڲ)��˟�u����]r�*�ibp��R���~��{Y�������E�]�)BB� �.0_?�#�՟�#��<��cſ��!	�+�0M)~&� �D,W�z��we��k����d��P֚�L��%��x+<
*�Eaj~� a}"�8m��P��ʉ�2{�FF1���3j�X���|,�:W�QF�S��W��05z���4m�"�Jt��ɴ �)�� ����Klq\8���?�*$�?�Q���|�&E�+�'��M���-r/"W5��B����Ʒ�y��뇅D�D�, �O���p'@o���7K�5��URO�74�"?�!�e�Y��o��]b+@�&�Mښ���M���ib�h�&eNݸ����Vd��M,#���ۏ��$�׮]���s�M�Ʃ��y�� h:>4����O���68���Z���	#6N='��F�YG)�[N����j��<�n\���&Q���ScFy ��_ueSyFx��9���篦.�lܪ|
���e�2��|V��)��W��+�8Y�f#�5�Kl�m��y�c��']~����Sٕ*+T6���~�ae��4�f��w橧�ݽ����Ūw�㳓k긁�3�M(�-#��y nd��[��J����sh�e���jC���đ��/M���[�M��q��DJә�ryR�Y���6�=�g���J6l�w_�����M���&{ �R��}�y�s?����dX��<��羐~����.���t�ͷf�Oە�Lp+
�m�����`�[9��.���t�d_:kSwz���D�U&��њ��l�t�����T�R�w��&��?����W����|65>��.M��2�t`��TnxG�%h9W߽fy�K���Pb;z��0%"�`����K��؉���8�\�1c�'�����$ų��`����4�(�"K��+�|	��e��RQ[O_և��ǂ>�2��א�IeG��+��'l��.�Ib(��4u��GS qJ���x4`�0[�ɟ�̧q[6���,���lD��Sd˳C˳S�5k6mM�`���ҝ������q���`���82����kWN�ѩZ����!��N��O�y��҅[�&<��I�����o����W�"۾�7������kM��w(�ضy�����������']�N��H�Ǘ�Mw�I?�������1y;��������������%ۙ�qLoxd6�5#q���t�бt�#vrI5�V���.8�#�h|^������asz��^����K-��$ztra��=G]"��֥u܀���z�����'t"~�X\�*J��&�swm@��1�xne��^���ko�;����{O�y�>S�\������M�����}�+�D:�NJØ�bB���!&#��4F1��ԭ���Ւ2�������Ci
f$�k���~�+=VҫJ]�o�q`�J!sB�
+�j�����;2i�3qD�Y%C38�-?AM�`���V�UI$���F��'���"V!��%*��2�1V圸��A�i�0�{�Q3��7���.��ݶ���S}�Sư�����ȑ!�+�	~W�.ZM!B�"?��
Ԋ�ۭ�q����2�����'�+��3R1�,�Z�_y%�7R~�!�NߒMw?�,��Mқ��cD_f����&��$� ���PDE�.�]ӗƆ��~��Y>�`�~�/6mX{�3��ԟlߺ����l�I'_�h�+���ō7l���ݗ���rn9�trvq��-5=\����<�~NC ᬠ鍭m��GY�c�k�x=�Ӳ�hL��+���$,*��^��Py�o{ʧiʸ���+��o�G��tha���m
�71[�-R�C#�������_��M)!�$M�	Օ�eC���^�?�,���Ѽ��_�J��]~xb����/G7��kA�8,MUi�.w������+�"�b ��W��y".��VNJ���}�I�ID"M��:��8�%��u޻gw����Էe[�٭w��~�0����^������S?'�P�J�؊9��WD),��ח~�������ig?<oj�f�Ͳ6�2^0D�ҹ;6#=����n���;�7��%i�Z8|oq�q�P������aFZ{�Q�]���M/�u�+�M9&�=p���w%�̆��T7V�Qd`1©�E�8ѻ�7^D�:��o�|��#���I�:{}��&��(܂���v��צ��G�F���&�[�����_7Ɯv������n@:f]\�[S��!�NGW�^��J�TB/�]��[0A�TAD��b�� R*& G(q��"���]��4?6�]v�Y�pK�돦?�?ߝ���/I�?�bt�Rz�^���c_L�c��h���GG�k_����'��>�j�`��O��c�O��>=�q�K�z��S_��է�qs]Z�~3W�܇M�����3�1Q�����[��6 �ir�h����D4�aD^��+��}�G�%�~�G?��t�ڶ|���2e۞������Rs�洈�vO�f�.��[�ݛ~��M�_�+���ޔ:س��Ã��/>���nΟ���>�Y
���dOԎt��υ��J���+<� ��g�K��g�>���}㜓�3��h~�%puKJ�{�˲'<�9醟_�>���L�k����b�΄�a������=��/�U1��?��K���'�����_�P8i��6���V��������x��\Pl�7(�"/
���a����6( �H,+>yUnŗ��2+�x(�x�U80��:��\�.� E&ε^�m�ф#��:���\�Nzl�vN.��ݹ�X�Uj�8&���d%c��^,*�Ŷ��C���镒���$��̷����g���VU�Τ��Oŕa~ʝ���w��2W)3�r.X�O�G�R�������[t�p�pz�8u4���|���:Č��S���0$ɪ�U�U���O�3O�Hp#ԉ&8ڂ��	�!��W�����\��|�l�g[�:U:�z�E���g��A�D������zl\�z���%E����v�~ӹg���3�~�������e�g�ȷl_<��}�O�b��_��M��{?���|�@W�#�o�j�Φ�#1����C6`/;�]�N��[�×�j���"]9��M��r��2���~�W��]��8���+�~���_��^��w�����^X�!��W�@	�iz3d��!�璋��޳���M���|(��8����Ǝ4���lzthCݑс��g�r��JеC�W���ϐ�y�j����"���;�k*8��M��E�Y0Kl�x�ȁ���qCjmm͛�:��6Nc�`ե������o�`v�;қ~���&�G:�Sl 1�5�@��ڗ<+�����N���uY�)�3��(f�a;�I��Sa��̬�~ ]E����_~ߑ���|w�����.|���0��R��糭�lS���~�u�fk�ccc�i��]�YZFY��������v6��*��R���5.�H�̌u��Y[;���L��`� ���|r�jh�u�tf�qD�-��#�L����!(�G�c� �I���,���85�"�J��og�WQ����_���N:{BHk` Q`Qt�ȸ+*:θ�
��:�aq�Aqt�Qq�A@�-BB��;����z����׷���9�T�uխ�S��SU�P�6�ÃؒS�$��u9^����6�A�Ը�;�՟�34]^�曐$L{�J`�+���#ݩ�-u+�!xb|��?�n�ͯ�U'��N]�B������/���=��3n^uq4�̛^u�I��؆z�I���}+޾�`Լ����>�Uո���bWQ��-��8�<V��K���M����+Usx�ￂ�����SO�A�q������w��g�>��ٹ%Z���U�-v�b�y�sT�k^�ҕr۱��'z��[�+�lӖ���+P
:�M2:My~t���4���ܩg^}��uO�����]mh��w�{��(��Vw��Z���'�ذ1Zz�
�g�^�o��蜳�r؝�sYŞt����Aw�HK�d~5Ȫx���'�t�O_�%����WG��X=���_����0L�&7=��)41':0$����m�uJ������v%y��eٺѐ|[<�%0_g�hj�X�m3)���Z��ґ���D��(}0�#v��t�4S3�0yb�J��͍J1J���69�P%���:�_�@B��A����H�6CC�1���Ѷ�o�t ~/2��q�0 ���^a?�!��?2z&b��L�,�vʈN�l��÷"�-|�/	� �Q����o_�&���2XD2-#>
��T��9�,�"bi��qě���'#��#��T'|��۪X��?����j�IP��T��B�'�9�0�ǒC�Q"*t�7ME?K�0��D]���[���=b�`��S���~�r��};��㝗]���]~�V��$#iw�W��j�}���7�=��Ol��N�7���퍣������"�kG�jPbY�GYМ��Y#����Cƴ��&��2sy�i|�/���8!<����O-H_di,ŌW*���Def�pcQ�}�^����'	Y@��/�����W�Y��Z6������U���ݺ�
-�]l�#M��.�M4�ic��IQ��r6�:�lŜ��N:y�=`� ��c0�v��=�.��e1/������r[��56��2��iE�[yR�;��O^�O0�cnɂF�ꗽԝ�⵮���#9~��c�����r�a��hR30s�*Pśqv�EO���R�Ln�p�����-O�@oҲ�_x��ϑ0'�P��Ⱥ�
��9�A�I�4Ԫg���;`0@0Se�QgW�+b�-cۈ��)����j�3����*+�Ur(\kz�*�W��t���)B��]o�����c�<��Ҍ��������lr/��qI1B�����o�����D���نStD��c#���S�ܴ�F���S���C�Rd�:ن����\�7|9��R���V��-F
@ft��ͭ)��PZ6�t���!�2�W\�B5���wF'��l�A�Q��cݯ�ϝ�җ���9��q�eYYT]S��?�{ץ�q�nԽ����^y�M�Ls.�-���¸n�	]o��h�X����~��!�H�y��>����]QüŮ�����9�YT�MH���0�=��d�v�
7�{oǬ9�mٵ�mߵӝy�� V�\� ��"��������z�cU�8G�Fmݼ�ǖm���P��[�����m����&oH-k����;�����GG�nFk=*080��|_O��S�o[���i��̓46����4�@Z�m"��\R%�CmA��t��'��x,�}�Q�l�Tt��$[����#FD4�NS��F	 5(��֚�.�9t��"g;_�<�̃�H�$���(+���c��m��(!�I�$T<1��3��s���M���n��ma��_ƾ�r��'J�#�%V�|���_I���w&���{.� v�@jFQߔ�����X%����ȔJ����֥mq���<����J��6�G��۷'�
@O��vUD�,{4Sk?�PmI���)<!��\*U5>�1M��b�EZXd5�0F�G�\�a7-3�n��h�������)a\���~`�Ͽ����%�-?��wL�D���
�e������h����|mt϶�2��o�v�v��I.ʲ���7��̲�.a���]Nr�7�Rf�ML����
�a�x
�`+��!�w��Sq�`���N�8��!�l~F3�V}�C]l=�������s��_s�C�}�ӹB	@gڳ!Q����|�������y�7;�fys�m-����b0���i�h�j��{�".�'C����3��7yM6$Y�5~�TҰ�Dr���g,�r����|�]��k�ܥ��OZ��1��a;p(�l�SB�qRu8��V�8��]'k2H��8��}���[7�6~�ygEo}�y��`SS~t��+�MOnӫ���_Y�;���G<��Ur��58��Q�AǺ'����QM5qyI��Ώ�G��/FoS��G,;���_���
lb����!W�������s�-������v�q���j��q��.D��{�� J-a`�*=̍���v7���i;�?�a����
=�}�V�:(��7ʋ�����6h�H6�j8\>��za^a\��_�)6����:�����mB�X�ـ��k��lI&�d��`�(j8��C��uq=<2��c�%�g�>w�����/]%}�\�w������\U �c��35D��w��\wG{�s�N��I�����^����0s棻j,�k�����&��vp������	��׈{�.g���[�L.�$i������+P)
c^c�Az]�d���u�MQ]S�V�ͣA[g6&వxэAn����n��������k���b?�ˀ<�������mٲ%>c�"�����,���	1�bS`�]�>ΨE�c�1*5��GG�����fT�V.�Do��LD�[;\��c\_q��`{��K�m��z.�0�Mz��Y��$H�p��4����ֈ*[dc�>B_��@kh�N��'M�F#C[�P~��M�u~L���@86�)�P�t,Y���~<-�����R����
&:�$��fy8K�0��~I,d��EF�|���d�<�x��B��L /G%��3��Rs�I�AhCӌ����~�eQ�s��>�<��J�m1x2!�Bg���$�	 ��$�Qp��{�Oy+,�?���l�;�~�T�C^��&VG-��Jk~�����W�~VT���[bϦ��bL�e
��p&�}i�(J�[U��oqع��,p�,���:#nŲ�c�@5� M����;���_��U߾����2�f�!�����g�Oǻh���?ܺ����~�h��y�����^n���8g�����O�( ��n<s��T'�f
on����3����������'	���;��҅0�!<������?��(n_���}��I�AQ�ήZ2���c��A���i��@����K����[7�ܽ������j:1c}�A%�l���PQY1J�&��
P����d�ob8I� O&V�0�9VyL�=mG�1K�����������t�_p��Ⱥ}���+��}�s�����G�-è�/q���������-`���΍�-Qɍ��ֽї���k�+w_p���iB׎ĩ�(��|,.4���?����j���8W��֖�^
�2U�:�����Y��������R6ؚ��)HE�T>�����;�z��`%���NZ���t�]���4׻��&�����N�9��m���r��$����P��W���b&�b`S4H���zM����EWǬ`<G�ND�H��#��%����H/������[�{��#��F��5q��P+���M�
O������d�F�Uc�e8�=8҃n�CѢ5�y�F��0o�@q�(b``� ���)��1���7�tk��G�M��#��i�����z��0�P����ٽ/:���葃ܐA3�����ȭ9qy�C�,"�_�v����hz����u'��_�Z�5���	4V}M%�WD�̌R���#��ޮ�s	h�S�e��u����V��)���0E:�]<�䪑3^���Z��	��j�[%0`Ük(���=�qL�ww?K/��п�ϯ՗��uw���3F9dT]�{������AO�"M�ZVQgP�0��n�b�X��G)jO��M�#H���D��W���Lb>�6I�#��Nè�	�fT��/g'�Amd��zf�qB���Gd��N+ l��dMmƤ�DFpd42 G0�-������GɱD�9����Cq4e�Ĉs�ک��`�0��'^k�̙|�G�c�����ٶ��Ut>�µ-�38Х�0��|�)"����hnSp��_�{!��+:��3���V���1E��6�$����]��Md�*UR�upڽ(II�=�C�ʇW��hQ1�K��@��k�X��O�@�}��Ien�E�l�a8lEQǴ����3}K�0	�Ϸ�[���?KA#Z�l��rWL���#ܦ�xP�qi3}�����Im{���?�ʕ���+Vt*�2*S��)�i��7�^���z��T9�8�u\���C�\�.9Xh���2��3X�k	]�Q6Y;�)hsq�8�nEy	���-L~�p}�)&�&�V��
��!�׎�ԑ�?F����;R9�n���p��	(��f���~���;��w>������9���-HG��5��(>]A��X�r9 j���Oڑ��լٚ�4����L����8Qʒ�������A��e+x7mw����{;�*]R���ʝ���&�\5�]y�nӣw�M�֙����ϋ����cV��*K'�[~���� F'��5U���;z8PpЁ�Ο⸠�1�l^�vKE���S=�:3$��<S���:�6�1���8����Ў��$c%e<�g��x~T����_�`�k����w���1y���˅c0�l�-k�C5@g����j�+�A@�@\SW��-ow?��ϑ�!=5� hl���I>�^�G��èp�	[��Ę-8$>��CD��dd8�G�3$�>4���F*�G3��I��C3r���a��m�2�p����Es�/��"��,�rb<��л���۸�i��;����N���W��k��t{$��&���aΘ����ˢ��\&�c��:��%�./�֭]k�c�,E[ 8������7������^󍨰�&nll�6ox�-[�HB�����B���s6kµ���̵�=q�RVt�v�s�؏��s_�BS�𙧶��(6�]�(C*���õul�R��C<D\_=��I7������\�$]!�	�8��U��F����~<����%�����í�ugF]=�Ɋ��z���" �i��y/�/�_��  @ IDAT�g\�"1��:�vz묿���3A�\P�#��P7��(4��`{Y��X��Ⳮ��KG<�h�I�Fb��%J�
.2f� �����b��m8�D���� G���>�h	 �L��&C�WeQt�%@A]�̝+�ԍ1HZw�܍H&���h����$�x<Y��Hљ�SD�Dt{�×х��6[r^�6�)�z��O6Ã�H�Z M�BWx�`Š�$mÓ����X��p/�3�B�h8&KS����8m-���\� &@ٿ1^�c�Q����݀�d�3�b̘m�l�h�%f�Ү�8#�Q8R���WnT�\�N�'�%y�
��m���h��g+R�"OKX�qP��;�w���o��k�<��ͨ}&e��e��w:Mڝ�o�����W�޹l��gm���1��6�mqˍsR(|FH��2IF�g�,�j�9�;�3����M�Z�5��Nk�F���aw:M�?;�q��� +˩q�/&�ˊy���l�����&"��ً�xt�qK���ȓ]u<��$�����&R$LB�F&�Ц5�g�\'LB� �T�����B�ͤ}�F���L�	��4�D�-v7|�F7�7(J�xf�k#��Ѭ][Q�>�ouW|�n��'�Z���D[��u�;�����[؎ɰ�7�A��h��)�hԶ	���:�����VH���c��G�dҌ11���ų�����6�q��n��y����`�ڙo9�Ao�ޅRf(:�Q0fgY���e%0�f�3֞�Ψc�3�EK#���=@|$��T��}�&�c�a7�<�s�F�Ǆ]4w!�E��AT���u�I���He�R�^���h����)�d�Q=�ph�7r���e+ت'y��\��D���G$i�r�3��k�
��5e�PwO�y�`��S4�G{�w���GP:�:���"������t�ş��*�`F�qǭ�����������s眽�-D������w��n��=nű+��[�߾�r��xc(�Z�������EF�aUɎ���Xwd]w���H�A���]��w��!�fA�o��e��6G�֬��١h��gtSD@9�u�?Pyׯov����}o?�&���f���N�{j�Oe�T���:�]��kј�?>�{'7#�-�HJ�c�{h�FWZ[�-_`t��W�{�o|�)�g���DMs�O���+���I����#����� FG]6����s�~(Ei� [�0I��B�n���(L��9/f�)��W�1��3��������R�i�\	�fQ��[�Y�������ȦQ�5�[_����fhwD&��!��cD�m�M�=~͸�B��cW��m�PQi4�������FzթI�_��o�\ N��8mkz�Ǚ-:!�̱�6)�AD�@ %�i[��ǣHٞ�)�gٞT}�s�?��t�� �,ˡrշ��n��}[ uE!X����#]�Z��N!�X�_j?��Xo�chq���3�2�&yd�-86�k��b�d6���<��xr�E��FZ�����/?%x��&���o5�p��+�,tI�B]�q}MItd�SO�ՙ'��n,�/�����W��(�s��8�p/~�����/�Xп���S֛pc�c�P |�eل0�\8��(x�����4�t��~m�Z�3�鞇�)+ss��Y)W��(MXB|����B��g)U���C�w<�~�G��}=�P(�Scf��֧T�D�t+�)� p��-*�L�싦˨�#��,������g/_�v�1�҉��w��۽ₗp�|�^G�qK�G�*��t\eo��xsLb�5\���5_p_��;����m�d5����׽���m�KJ�;��z����90R�6!6 8�ܖ[��E��~`�FQ�r̙c%c(����3���i|��/��F��吨�e9�"�\�DB8�{=�H�xX��w}��r�XP���p�r�O�'����+��?w%���
4�?<��}�[7��ƹq���PG<������6jD�ި��,��3Ut,�Q�����ٱ��Sn���rs�2V`4�p5�����r�D�����notxAUcC���[�2��Pbw��V���;�����箼�{�|]�ws�^q����qIEc����a�)Y͙Clm��z���׾}��r��ܯn�������~_���㓎[=�����oxu��W�XE��@t��E����r��A��Y0Z�n$j���>���I����;��(j8"Ϲf���SO��ڴ)\_�<�m��h#�͢����}��v����}�c�崂�:��Q6�m8���q!{�@C�����:�p������	w��ᠹ�<�[��~�jW����M7�(o>ʾ�k_�L��?���ۿ�0��������Q}}�v���6ގ���yuq�. :p#��� *z:�т���0腜������r��k��uc�rm>��i��_霆������[��l�S̑�}�U�f��X[ <���'����R�P����|2h��`,�|�Y0*?a���UK�t�0�B��Ӕ'���9�U��	��pc����h�#?�6 :r��U6n�NX7����D�a�(+c�6I��'�򑲍��l�=zl_����?1�^��7I|��Ựe�f'~1`"�\(?��?�1�j�Z-Z�8K�o�,<̏�	*c8�e�菅�H�<I�cp#Fn���P���m��$����I"���2�$������5��<ǥ�H����s������8tXZ=p��/~��O*��UK(�����f~���q�杤Ϯ����·=��9w�܇Raސ�c�H���������F��~ePSy	y���2��4!N�i��������}�Q�!����P;��\����u��������.����Wn�8i"g�DN��7t�?����/�;��v�q8����`�Ǧ�7A�
\ا�h���Ǘ�~'#R�$�y}����F�u|������;�AuN���(����Mc-��Q�H��"�<[�j��t�H+U�CO�u1� �X�se^{�.OJ�8Jk��/o��mܴ-~���q��́��H�JZHx��nq�x�+��jH&4
*�����WZ�pxxt�ZCܕ��Q�,уF���䦴}� s^!˔<n�M�D%�}n��@���p���F<�W�e��vw���ot'�p�[�z�����m�_�������]ϫ��*&�X��>5J���s��Mn��nW�����ӵ����7��*��&++��P�4�֛�A��Rq	��l阼�U#�M���l?���.@Q�S#6f��	�&�*������#�>rϯ�7�;�H�>i?�W~�w���8��я,z�E��`m��G�j�Y�����8;t���r$Fu��a*�bQ#B�6��r�V���Í>��B"���,���P�`�nFt7�-�-ҙ��^��&�$�C�m��/|M�O�:�a}��ϸ�N�J��;n��/�w���/�];��jnĝ
�u���f��Bl�uІPK`4"X����k�ݗ��F�q������U����x�k�)���&bn/F--=n.Z$�l��8<�������^���K/uu0U�Y$�0�ϴ��"���6f\�TO,H�z���9�	Z��TL��7B�9�'�	Ci��;g�~�s�l�F�V��N�f����8�*}[��W�b����L��,���5�j� �lSK|�W�b˭C�::!#$!�
N>�o���S3�pȄ�!<�{Yf�}����ϐ���Oq]J�I0�rH�+�_H"�H�����^e���cpA�2�IR�O�x�E�d�\�Kҗ6
�GC��#����g@G��lK�d�,l��.Ʉ0�H��Q-|Z��Q�Y��� cq��In���:���O�yܒ���W<��_:����	����O8�2���W����?��o��>�Yx4≬O�0�r{�z�{������4�/�"^��n����h��i���~fS�2Z���q%��k���ѱ1�*���s>��l�����v�4lGͩ��9t�m�\�b��IE#���fT;H�hj�$�Yv��ǻ��i��;��^W欮P�M�*fI�λ7���+*B�s!���2Q�}��x�Uj�8��z&Mp��H��w����}������7�t�x�r�ܹ7^���m�lb�cDy%n�ٸ�=�b=>:9̠�e2��}[���� }P�0	��:ˈ2})���9jAyr��w��������Ք�E?��WT=ǽb�¨yނ��e�ѱ����Y:ھ����5�v[v�iZ����s"�Y��#�~16�З��l��wq���kx�k�.�p�o^aqi^1��l�Nb�`�V��3J 5ojc�y̏~ S��"��8��O�;y3�v[����PTRZ��}N��A6��=�;�4�b#Cv��z�)����}�g?�Q�����~h�>�^5�0��u�l���	����F܌��誽n���F7̩ԘpF_��䕟�f�#�?���]�����M���N�dg"]ӿ�����o�K�|�|w�g>�ʪ]t�[��U�6��"�����賨�8��j{�FEޅ.�O}�:w����%�^����]�D	������C0ڙ�2^��9��Qo�}���p�?��͏�*�z����CW}íX4��k�q���vCc�S��?n�=��n��^#��z�Q~z��!�U�1u5?�Dq5���֣~��ȟ,����A�J�x��&9+�ܰ��Tc���s0˖�d�N�'#ZD�W�3T��_J@��Y�i6Ah#��I��/�xM�M�U�Dl�Sc��i�ф���;C"�P
~	�H�8B[�ApCB	���4E ��e���I���KѤ���(���L`'�d+��Ws���[Q(H�Џp�����V��L`&����3yCE�j,<I�l�:��\z�hҿ�E���LcR[�&L�p|��p)@_*jY�)�
1���L�e�b�$�oN�U�-1��ne%t��FC0���jt2���O�ߘ2 &̑R'd� (�c�GYYe�̓H����c�N^�����(>��g��o�	���t���t��%5Q�ܵ~���9e�M�:��B$�SRl��V�9���.~�y�|�iVܙ�)�̧m����[��U�:�2]�%Z������V�@|����x�,E�1�p`D:=�4����h��OZ�Lh�3m��4��;4f>�� *8c�����}nyM��튫9:��ri��p�wm�l"1�E<��R�"K*\��67����!���c���G/zы8�<*V+�y���}�v��}&�$�Ǎ���R�������$�����#�]m-J�
J��8i�=�s�l���u�ə}+n�)�I:Z�I�x���FmD��CYǗ��mh�G��*׹,�n��pg�uV�^��G+����۰q���~�J*��Y/>�u���_�����s�@�� ��+��6.��Yn�U7�\��9t(����&���;��z�֫�R�m�B�>�&J�U�i8T���:��XR�[$su(�0+\���²��WA��tY����}wϯ)��V'�EYdc}��ޣY��,E���*w��I)��3]�%e�8�<�J�t�+�y;��}�����v7Ŋ\II&no9��
���2��1<;5�PmGK[^{��0�ͻ�Nn*>��[�|���@?c7�k��ǟD�I��;]u�5�����C���1Y�7�:Pw������5�ǯpMp�5u��D���Sn�/�'їW��+EI(��y�)�'�����u#~:��3�6n��ڱ��z�y��U�i��*�;[�ܒUkܮ�{����G{ܽ��Eu5�������=��[�d�mO��g�����p�1K�j�k�}��;*��s���vp?����q�YIyi���V��po�4M�3=bF}�ɘK�q�V�����kl3E��Cw��e�g
� ���� {L��q���T�����9,�xxڥȟ�QI���C��ns7�|�,!쒢'㏘F���P}�'���y�p˳�1tS�8OX�;�_�X�[�o�4�i�4�R��VFO�/b�&�9�!�Ύ?�AR��68��A�-��@�����%Ԩ��8�ۘ+3�K�D�
<ߌ?I� Г����`�l�W	|�Be�+�����iG�U,-�<~�7�x�
]�1]�E ��,7s9Z�*g��_���k�S���1`��	4(��i;�����8�{`㮃�㓽eECM����!sΨ�t�9�8Ψ�,z�����4�!/�������]��-!*(���x��Me�atp�����������r��u6t��S������K����������3G^w4S����#.[Z��,_i'jy�Z h���L�G���I#�T3�糪(f���VW/�x�`�?����ZH`jy��>���x�Ms��w�jY� �`���M׼8_.}A��4�H�t�@��r&�Ɔ���]����z��=�V�F�����&�(�L��f�(���1�$ E��%ގm:eIԀ��ߥ�3d��3X>�>_n�S�j��b$e�ˌ�&�^&S}�1�ee�qC�a�K*��l�I����0Z�$�y0e b���"**.��Ɛv�s
}=�$���G�4:4�m����/�s���S���bO#���ʹ�J�#�L[7���q
/��*��^I�%6�F	���/xQ@�"ތC�${𜙢g�b�bڒ^��P!,�!TAc_u'�ڦQ��~nR�JRZZj�����R�	.Ԗ��&�\`���$�x܏�݆��q�p��B�Wf&�޶n��9�?��]y���z����t4�᰾�gj
�����]?�Wńn�p�P��Ky���m�_7�ʬ���ҥK�Ѷ˧�D{{;�Q�I�$��v Z~&�k�\�f�G)�N���S�'5O��Ctt�І=g .�OrRj�QI5���3�o3s�ǘmi��*���R�*p�SA�B���\I��L�ąT6mB|�@k�!b����I:�����럔�M�x�2�%֒�;ry�5���}�\֯�7��������G7��񺗬���H~R��}���C��N�G�zxcx|ܩ�c�O|�8�q�)LV�L؉���$Eɸe���R�4��|M+�ܐ�'"VR4�2H���&��|&�[���K�6�&n�m`O&�YV9��,T����'0x��n}��
�D���¼���S_U$�$@�%��ƽ\�<_ܐJ����;�q��<���M����������7��cݭ�n|p������*�/�k�/�f^E�L?ы�_$�3q	?* 8��D84��
�WQ~
�
��7oݲ����+�-dB଄���ϓ�ip��"a)��p5��jTk&T�gM�j�U��$ �Q��:-�x���ht-�Ȕ�m�؜7��)A�(<��,�9G��/E�k��2���gl�U#��'*��R�r�L�P&��+�ɆRI�l.00)1�2���B�/�A����T�4�jBՄ�#L��������c���3�"f>b���AG��0j����lU�����O���"���n�L䟒����^���:�R��
1fh|��K�!z��I׵��b��^�"J�QO�V[V� �D���q�f�$�REf����_l�[V�ԉ��'�-���/L�V�bz�؊�y��|D��	HGݴ$���<�s%ĹY�&%ޡ( YnҴ22�Q���x����3:��GB�0��QV��1��%�zc�!��^������P_������ْ����!�pQ���ቨ}F�s�Fܒ�]?g�z���sC*;�&"ɚ�?�u�ZBҲ
�X�&�m[��r��������&Wנ�����m6΃]�(���?���<IT���e/
7��iW�h��L��E:�E�;��������T�Z�묊���a��iѭi��9y��i�:>��S�����Y�!��\ �:ES�Ǧ<)c��V��QJ�1�Ù§�'�b�,q>)�H��ۑ��� �|Sָ}�i������E:Q�J�����c�=֘�D/��UM,�,*��D��������?�6��n (���f��JK� s5�G%J_"Kت{�h���<+q��=B��+��6F���a+K�8>�4�	�����x*ҩ�Y:�S�FD���E�x��t�[8U![�6�7M�S���E������0UN����X�"X��e{|�i��#@0�
������9�r)Gi�v���o�UȢ�H}�ǰM��r�2nb���JN��"�;Г��_��l�3cC���mQ�8���?n{�V�^vjڵc�1�9��:�<�I
�����ⅰt�������P�S>O鄫�42� }�2`h�9�!��5Pu�R����(�%���$� ����8c�h>�W9�7����q�X/�39283�v��N:�L��0y!*��GƐ$11��?0�qrZ��u�]������B��BT���(猄��^��X��c\���1R�`��h-_�b���M)c0�Ε�Z��U�����0�ϡj� ��3
��g��##Q���4����J/��idd���xք=�I�-����Ó#l+I�U���� �:.D�
.0��&����-KOj�U��suf�4�*G�2�^=&z��ф��2E�!��nt��>�����|\[��Y����	v FMaf5�V���v�\�t/��	�~C0��')/��]~�5�A�)+��m�h8��MAy����pg��<�g�Sye|�KN�7�0�4���W�t���Wo��{l�NW�0~�T���z51hR�ȫ�0��u���1�zG�n�A����j�i�ʐ ��pI�Laa1���`��oPB9JZ����fI1
��.*�V��!�؇�k��c�VNIɯ�r�K�L>�9Ɛ��?T�gF����!x�¼�
w2iA��,��O`��y|�����֔���ae���+�Kb�"[�ɑ��$�?�Dn`�ļ�	(�*_N��cH�FElB��?�a��6���GmM����-�
5<�<����*>��S�3�� g,���{�j��o���9� L�/@����>��{�C�e�aʎ���÷���?.|��YD���#g.�O���$>>qMy��Z���YJHE	@�����oh�$A&�2�,�?��Ğ�-fW���%����C��y���/i�Q��X�����l ���PfK�N˅�J�T�"�.��K����,�Ȍq�b���!�3�M:�<`Y9���?�/�3�ѫ��#��g՛W]���4��?в�PK�"
dq>wʈ@}{*�ٮP�!d�4��tOO�����k��C��>��+Q��D��.��F�}c	p�cm3�.s+@?�yZ�I��=�5d+���R�,-	��l���N��+�����X3�j"C;$ۂ�C7SǐT%��)I	��l1&�G��ϐ���^��6"�G�Y���	���gr"\�q�%�������g��'7. A��0��6<�+>��"���C�#ZPabkm�J^�Y�h3S��3�3���@g�Bx�&Ɍ�_\�CQ��b]�6SB3�<�Ro��q�O��6���+:D�e�'0� E[��`���@��6�&$�>i��=���1TK�	�(J�H ���z��d���W�d5� =EpaĉIJ��:��b��y�00��j�3::7�6j]l>��I#i��Ezn$m� =��h�>�$)v\�e)۪�Z?��^�!ԋ�ڹ�F$�q��㞁F��z��Fw��in���d��b^`�����<$�S��JPL}��<������<��$�D����'��D'a�3%�� o���X[%?
��@�$��P� Y�94&+�vs^ml�*�~ E*:������DzU��1j$T��A�|�_�9��z� baK���jcf�2��[�1�W�$�$��@ߖ}.�-`����#��L�"��0��%��q�j����_p�T�qd���tԩ�nˡ ��W۴��>M�y� øA q|a�e�'<1�n��-�>��c_������)�Ъf僬��9��0��kZ�O�4)��?F��S� ,�o
���pky
��[��P�r�@
�R���`��r&՝�?Z��_�%�G���emբ Fk(�X}P�����e�7)i�1� 8��t�b"�F<��<Q�76>�W��œ���aB������0C�������75Q:��4捹��3�Q���ak�ߊ��`��s��Τ-�;������g�(L|zj�k��u�y��v����C�����Oy��޺���=3#3�C<e(�;���m�v-�n*�q=�l�
�	И՞=��vÏ�$�f���0j����P,L�&bk���_9�\�G�8bR ����e�ql�1q���W��fBǃ�(3��J)�%�6Ak�kJ��|C�"8��')M�0�0\�aQ: �p*��Y��/r�N���-��}>�m�|�����Y�N�0�����8���P�I��5&$� ��`�Tt{ȍ�'���f�s6ʳ��	iKڦ�?R($o	ʨr�����F2O�U��O�`��s�t�Dy���<�3�$kT]����W^�V����|R%pyI�d²�3)�ڕ��HU9�$���L �\���h+�׀�x��6N,
��$bkc<d��t���S�����<-X�I7��D�X�,0�,yI������W��D�Bgw�g�V��� F��8Z���aW�V./�q� �u�V��^r���N5L[�	7do�Y�Bm��)�f���b2���1I'�L�@,����MQ����yBH�[����r�"�66������D��d@eK��([�0�0�?�e��EZ�6|�Ą������~\�VZ�����W��
oD4Um�DJ����g��1�>�Z����{�� !�!Y\-P��K h�J.s'��QAǢ����6��>�����Yz�leVq����t3����/[ �|��5�P~>_�JB�/���Q^���,�n�P��m��|�|ƒ�RR�f�Ga$� ���V(�$�\s8��<<��^�{ ���փ3��e
�OT��Qv+Xlp�9;�*��*`��_4g�.�4���:-�|��پCJ�	q��0��8����5��=��i~e��nDv̓�k|Ւ�����hM��NaҰf��H��S���g���8�n���i�����0�j`F�n6n��qxyyU>�r,ܸy�Y���y�' �=3#3�g�;[`��[���m/��h������d�����4���S��A�Q,�&�}�_@��L� s�Җ�;��0f��
�<�Ot�
 *��=��{B�?5,�1@#<�1�jw�&�2���fI$�hV��e;*�Fǁl�BP��)�0�k����F
M0ZtЉ�P"�>�ԢU���*E������� �t��j����+�AL?z��d�@�ɗp�!>�'H�2�M�T���1��G1l�ha��ާt���;)�RC�-�T��%[d(�����̑��yސ���j%(�T]|�@��4�b@C�I�$���9Z���?F�f����L\���,���ܒG�&̠QM� J� @4�*��Q"���_�m�TMU�$<�n��g'�d�S�+� �8^=�P��f����ۣ"���Aʾth�FCT��c��
�ʣ)���|!�V����h���Ag��_aA����"TI薟� @Z*=4v`��RΌ��Rs�VtJPJ���)ծ�SA�
���!���Ym�#��<���6з��B�08��i�6JR.�RFU8_�l��
K5�m�o*}�O�v0>a(�<�m���Om%ߚ�RyZNp�5���U�S��r_&,��h��q\y�����F0���5F�W��?1Cf�6\�g����̪x��Z���e>��A}LHl�PG�( C��B�����i�g��)�_�t��"LÛ����g��x�b$	�>k$� OK/�Dǲµ3��g��� ���u�N�Y��CI���ic�Z\�����I���a����)�;w5��p(:�8m�K ��[0C�~�
i�/�����5}�g4��`����X$�u��¢qT:�;�ό������[���Ƒv+��o�Ʉ�r?W��;��pG��xɞ9��ĸ��A�f�M�՗:p����W4�mꏻ�Ǣ�)%RH .;�;��0�e�m=����s��OC�pwo\�^H�6�"Y�v��I*�� �b`�'�=f��F�4��7�΢B]o�u�����i�cJ�:ֶt� �<�c�n�#��`�%��g��c�+`R��vf��x��a뀧:$�B]1�tP
y�m5�A��	=S�2�I�2��tV��&��+��6C.!��B�U�DIᇲ�z�D�D��1I����'���6Q�
���Py1�3�2��Z�-:<����ڨ!�$�D�(O��w|��-�'�1F�|��`4O�m���T�ja�1a���� Y�h�E��]�bQ�d���;A��.��{�%t�)���f1%OP�!�1Q&�I�eT����&'�E��t�</�6�dlq����E�8]RP��e8�j^�y�����<��(5J9u֩�N��f���yoI܈$�?�dH�c�����Ǟ!�U�����\e�t0+"^u�@	�C����X��N��<R����Y��,	���`!��$�yb���YuE���uX<K�P�A����l��0����@�1阿T�%ш*�aJ.�|"}J���`+�_��8�w��ڈ���!&�6��M�+�8��ƧQc��TP�~���Z:�|2�&9!��l�O�S�'��,�Ri�IX`�Xli5�������/1I�9-�� nN8�0������۔�T�ϔ�t��%1�ϣ�Lh��+�%e�X�&���u��D�2���.+U��pe�ʄ�����#�_�r58��>ԩ��(�v���~����Qt�!��
&|���@Z�;m+���RM�K�qõ�����ݯ������p�D�*Rd�2�1q!�b��� '�ހ+�I����B��-;��?�
O��-�Ӧ�B�`�TS��w�%[qC�`g�t��:��=С֡�x?T.��p����--sv9|�������GU#�IܝF��D0���$o8��7���4��ɂ�������\zXٚ�:�l�:��i M�;�e�w�� ��:1�[r�(�BhQS�yR0��x�x���5$�g�A�#Ӗ�J�%��������#8	^k�BC�߱5@A�������� -�T��ˋ�#��L:��y�p�G�sL4F�*ޤ1"�	�h��`�2>�L!zb5ª��|!@�9�_�i4�'��/�B���31~�$	�hr��v��I0V~���S�fÜ����I�cW&�)dE��_��Əf��H_!6D��)�����w�i����Q���F��wX��r���Ӗ������U	����$���-��55+m*C�1q��TH(��Xb���e%y&�
]���_q��?XL8���KUm�U� V�2�
��a���R	g�ts0���a��#�4�<�ҁtb"#����<��л���]�H
��(W$X�����@mf�v[X�+�7�c9��4��(��6��9���&Q�meHI*������an�N�T��Z1WC�2�E�͛�����Vչ�JT�"me��s]ň�ئc��D�&5G#��mML�
�j.��L��1��1��,j
����O6X���s*��iT�(%K*���(e�	��Np���U�S�^չ58kT�ų8��3ĵ�(X�ėa�����`�+�
�-���ؒ%|x�ә�C�����0@:k'��s�4�B6F�H��xiXi�"���Y�T�$�����F>5f�_`"A1X���2IX�mF�G�*E�l,J�P�K~����Kh<�$��T��Dl��\�re5U�� jh&FF�Ҽ��C����'����/$PZ>��H�;q��BX:Mڭ�2��s癬bV56��lxr��{��e�-�p�D��w���ӄ���������;m�������o�8�;�!n��/������_�C<��0�sV�ކ�<�]��h�i��΋�ʪ���������{�u���MSG�M 9��^�D�/m�-CzZn��H��}�.;�䳆�ʗ���VF�u���Ga��˫X�*�o�L,�	b�h�dÖkI{N�	̍o����K���=�@}�����9u��pET�IXi��޿��v���>���D��g�8/�w�߸�;����{��zw�};�Ov���\u:���^�|5�r�]���j��P�4Loo���~���.F�P���h����J�]��[N���|a�w
�/�-�d��	Ŷ����`��xy�Xʃ ���ɣ�l!�����-B�y'�&NP����.����F����F����},���B=m;ť�b�QhtɌј����B��(��%��J��K��#�|�I�B�$%��m�)_Z��r9�6�l}[��YTK6fH�Z�D�?�X�(�՛$-���������B+��@�e7�iӦi!�O�����XݰԤ@i®<ib'����Ôh"ǨjD
�����pa+f�#���E����8̭ͫF��S���္h���ʊN)��/��5gC'[�D/�J�
��C��7�����SOvw��7qKWV8��l�2��a���P�0�D[��JPϠ�l	:��U�2�~���@d��'i�W��>�Eժ�G� ��:Bb�]��X̦ha� D�"I��z���}j
�Պ�<9�� ��_(F#�'�y�J�ˏ-N|suAAAW*��	����~�Q�*TO�I�Y�wR����6&G(��-�`&���9"�c�Ï#	��4���*��T�Tc�!��&�r��(9C�]RQ,�'0���Û\�J�&!j5<-mHi���,�	��[�gh�:�������d�1�4i$?SY���w��{{A]c��I�n@!� �tS�#9��`�m�9�{wÛ����]��76hieFb��628<�*��TY<2>2�`yڜ`	ǟ�_i�4>�[��+L�)����r7<�e;����H�x�V��m9��N8mm���n��6�ߺ���_���7^v��UǮ�TRR��@��+M��L�Ca��u���;w\{��_?����Y������GKk�7�9�"���bF��D}\�ѠDGH~ࢰ��{b����&ϗ���ЧX��8d�!;�x��h�<�_ T�ٶ,��:wmvK�\璛�3ќ�9�5/9ͽ���%���9�=�@9�*-���������u���s��m��Gǚ��;��@2�G��;��:U7Ùs�_��#�D��dj���@�_/iX��'��	a��W��4���հ��,K4���/�7��#�ā��0���Д��j�ԪrMI�$U�e�K�A5F�o�!���j/LBL�K4�6���"���DV�G�"�h������= E =�ŗ4�*��O��Θ:*�%�ҴG�5<��M��M��fT+���!���S0�ja�=j�$OjYy��',ipa�e�N�����X^��j�h��������B�L}�a�+I#_�q��r�����(g�e�Mt1dz������ٽ%������b'���/�@�]�.��?�w�G�5��2�/��1�0p$el�r(Lh˄�l�D���s���n�b�0ƑT��ݫ�|�Y�a�-��b��e2�v��a���͐Z;�e#��m����(���c��`�(nv⟤7&`a�b=�[Ɂ�
K �C1_�
J�˓o����9,�2�f���r��-޴�Ϛ�f�,�9��@O���_�jL���И#��Q�F�*04��?�����g�Q<�x��`jڲ��8jgVN�c�\��B����ɬ�CQ!*T��S{�6�o��worO����ʆt-{��L�;�?�N��݊�6J�wŧ
�*WV͝[��W$�y�Бv�0gy�9�(  @ IDATmkZ���	�%�zf��s��	Sa�O����/?��/w:,�VXڤ�����H��4��c�˔�k���7䎲����W�~��755u�����7��77~��w>�k�[����Ѵ�l�wYj�N�fI�EYֲ����~��[��g���MK�=���g�����.���?���-=��4�s�B�6�$�������~:����0�,2sn�:�Z�j�o�s((������n��h��_��lo����]Y2�\w�?G��]��o��=��8�A�A� @�x^Ct��3n��E�]�� J�������n�w�5�����D�67D�<s22����R�ԫ�[C��⿚�jB���c�\�d��Ռ�S���X�oS�.2?�Aq���`�G� �ҏ���8��t~�q�Ђ�@R٢M���v�Y�D�@���A����#��Eaj��'v���G�i��Ot&߲CX�0�����؆Cvp��TvVn8�m��A��
ܔ��I����'��-@W��s1!H- K�0񃒆7DS~�F3��(��G;�H��%%�n�S��Gzա}���R���3ɏ�O�����%&�5�^`C�5���8�M9A�CEK����:?�j:�/y�~�nL�����*ϪC���ge��'4[�����x���W+{�j����_����t��DU��^����7����0ڐ����r���\��9�mn�2Y�B�p�28y��u�i�f6L����G ���O��1r*Sˏϓ�?�{_�jK��lk[�^(����-�M�E�Ў|�\x���}��/�����g�N�Au�Et��,����c�����c��<=�h��IW�Xi�d���g�f�^�}3�2L���M�`,փ�Z�ӍWa���������L�8?�������0�҅q�������J������� ��Ri���2e�ku�v��UW��4n�R���I��C�'���8���zbgK�F{�>����~Β���7��=��V�i�ӏfgFn���)�Kb�[�Ls����/����;����/��f��]lll�}U.��A�_�7�Eb�Q�'���O��!�[4����i�7����=Ӥ�w���&3�A1�A�R�s��h�� G�2��OlqN_�^�k���O���P�=9��M��l۳o���KO;�[N=y�f�68�`b|<;2^TV4�訷"
���;�{�<�}���<����w�qk�ZܸlE�����K,����'xkj���U��0��
��ӹZ6�����vB��^�F/C���t�̟?�	�a�����G�����n��.w���;x���� �:�Ɔyݞ6����6m��֜v�;��e�?Q�2��JyxIP��pU����������u��H���/�$.�\>+�|NfH��n���1;��!�>F��!�1mj���:Io4��CȊ�Q�W��@����1�?�ա�1�3��8�P6�� h%$�VB��1�y����P��i�k�ڀnxT�xYl�h���(���z�p�����eq5wY�r`��P�l�hS��}5)����9�R�jB`=�[����Uv�H��ӫ	C��XX�c�%�r�Qf�A�"�j��D�k��[�EW������ +eE�04!Z�C�l��Q����ɄM�*7B��	o'� $�I�k��z�HҴ!�2D�B0�JL�p�����J�b�\�B�
E/7�T� )k����x$;ՕW��o�E|��'�K/9�n#r=#
d���v�� _+kJ�I����S�Q8�y�IH��^�*��4b(�x[(��M:Q *ѯa�D�ȷ�-o_�槢�E߳���S��)�n�6��5��R�T6�4���-�Թ�>�\|��7��E�� �T�pb<��
�	5���a�" * �jP(�O�*W�*|Z�œ��W�uT��K]fAE�I ��}_��& R�\k�¯��+O�Wn�_-@P�x�o�/�M���/M���|^�ց�K<*�����&E �!A����CJ��<�d��B�xy�0��8��b��2Eq��d<�u��^�}�;���޼m뫮�����{��/��@��OT�f�����۹s�����Ӻ�U/��%y5�l�-�C�m����#����}�ӏ��:S^� ����=��I{��;��liB<���!���L�tjZ+�"93�c�U�=���L ��tw<�ɝ�C�/~ͥnýw�`�[�bEA롃���_#�VV�eO��̮ޮ�α��:^�.,(����wV�ֶ���6,h�>��ue#�Ż�󆫛�����޾ߕ6.�JdU47���s��4y ��S��Ĥh8�oznH��K�� ��+LqSƚ��B�F�����@�>w�g�W�f�E�k�1'W,]�栻�7GEus�~��_�M��yx���؜F�u��662�20�� ������ ��6<����5:��&���Sܣ�=ej�y����H۳8&���;���ʏΧ�d(W&5$���@���X����E���<|G3̣R�k��z��b u���	%�`�(M-��)}t�&��>��a#&��R�AF?�ՀcTkբJ2�I~T�Y#�W *'���
J�)HŅ-(��7)��\����R���Jb�UE�mt�eF�������i&�����E:�n>�7%L�?�RV&���k��
1�U#+c4R�6�i[(�ZO0E`���S��VFS��/��T�%e*���[`���	�g ��@����\���l�HT]3ǵ�/�m�ۇ6��GZ]o�Q[9�9v���]�����_�&��nS^T�Ėd�Τ�����m2Wd\U��A�$�V�"����O������ʲ��������Kp�GGY���m�(�	˞�U�_���%��s�Ԓ�M��,hU �Ne�Y1	O��mi��k�'��^$�JV���p����)��jd*��ʣ!��P��Y- �x�o�|��ho*+CU`�웈ؔ��/�?ÖoתG���&�>����zH�#J���[��, F�O�.�k�!c���J�5�W<}�3,&�B�*���>�d���SnU{>,ո^�� fcS�Q���La�q�����O}���w�������{�^�=�m�H�f�?�����A��Í����~���?����P�x�^Ў�ˢ���琲�J��x0KY�j~b�H��i .���$�$��#�?�7���T��f&�4��a3��g��"a\�*5G�-�a�`���(�w��X�N:�7�q��ھ���_��33�UU�����{��y������qn��BoTR^�?QVQp�)k]QM�����
��+�������G�`��Q9�(Ԣ���O�q���"kCFU��M��p�X|˛��[R�˪v}<�0�3�~��_���5��UKܗ���h����;�.޼�5w����vw��a���L�r��6�"=��������{xy}�;�r�m��t|��Mщ'�ׯ��Ӽ;�;���FD�b��&1}h@��&����vJ.����eCq��mÐ���0�ol|��mP:FS�HR���fD�gńH�`%���(�"H�D]����{&�V�$��4�X2��[|dl�Փ˳��I���`$[��aIbk�W���T�vQ�4L�̔�$��b�(�b��������l���������C�+�d��a�o��CԉnFYo�?i�V����h�L�/Y��a�DA��Smj��]���V�Iy�=�UzM����e�o76lN~��GB�P��M��
�h&n�p��'p҈VI]�I ��T�o@�r���$��m��u���v���Ȓ�e�j,E�����&G��q�MY#��a)��-�W�8�$q�Ж�)\3dYK���L��X�[�/1����ࡶ��J�Ky4�L-D��|?��_og��ir����{����{<Kz<{;�cc��d#��  �!B ~!������"�0�(Ax�X&�&ĉ��1vb�سzfzz���}�����V��o_oaQ����TթsN�:ujy�r�5����i�S�
,u@.�N�Z��If�JI���L8�C�ƚ��N�lP���g�$�0�iy67��V*�
4F\S㖲��[~�%�©�:8�	��b�����ImP�±5B�p��7]�P�|�7Fم�j�Ct���BR�N�)�$'<�t����~��v��:U(�6~K�<�b��g�
��L��kO�����|n�m`�{C�� xLȯ����������?�۟9�3�����G?�����?��/<�裏�-l[-�2� �� ?|���KO=��G��O���o����}��˯���}�G�~�|���t����u���纕��L����h�^l/V�f�9�:��ĳ�[��џL�������o�'�'Ó8��L���l������[Z�&�Nѻ��]��G\�_f� ��?��K�퍛�c����?Э?���i�hkx���(��w<ѝc���K��nm�.��-\�xq�^.����6�;���o�����{�}u8Z�Y��jT*bzXX`���{����Y=�6���!)�ƭ����ٙ�u�6 �N����(?W�̭����������[��������4�W���rw|��m+,s�nyiz`oi?;�'|�áv�|�g�6H�r�զ�N1������nv'�k���Kt�;�#���ݸ�[�ҾJ����>p<�����Ph���M��u���*p6�i7�ГC�ɷ�
�l���,к�&萨�ɪ�� ki�!	��Ȁ X�E��4@�=Q�=3j����> ���p�/��op(�� MjT�4pF��c�P�����3�릔%R
���T�>��^J�'Z"�Q?\�b)k"�%��8�pKv����N�k��rP9�^62w������A�R���{}!P��
��Ɂ��-��K rɠ�����X����<��7g�����R�0�;9J���8�m�R7�t������]�Z���>A<as�!h�9i��������9_"���q�Y�TA�U%��X��pLT�=��
.uf��+x��v-�,�xPQj�'�3��`'�br�O3�n����2j�0\����zxI�'���Z�oݥ�Z����Z���i��y"P-��u�Y���y�����\'��l�\e����-II�]BuɇP��E�(�
/?>A;8~��Jw?��S�_�M�|��O��������P�����t,�J��x`�͠�IKW!s=_��L�u�~�Y73����\W�ڽz�����'~���O>���'�?�����������o�������������^��'>�y�ʃ�l�[[[�|���}�ӟ^���_}������������7�x�ʹso99>��E����O�W���_�8}~�x��W�w��2\��%N��fz~�-N_c�铏�F��j�aQt���p�C&�c�v6��g~����$X�iqg�-�Yzg�-���pM��;C8�C�Np�r*T��2LJ������۷�����~��N���ׯ_����'��O����P���͛4�������h�����n��j��#.�����/��b��+W��ݽa����qbp6��>��Q9�M��g�m��dR��s�B���N��>���������j?�z���5767���W9/���Y����/�m��/sa�k�~�֒��'H��B��rp�����%^�ͯ�t����t����ݻ��޴��^|�A�h�����pL���6�k�v��*F������%�R��I��˛����:����]Ш8:[y(��A���俺��+ˉ����f���:܄��!�.�ɸ�CP��0�d��	<ɥ�gF*6�q�^�x&���j�g;�á�+F;7]k�v�DK4ݘ3?Mn-�}c8�}Y ���� �|V�J����R�W`�ug8yM�i<�??�&���yQ[�9v�Y&LZ|b�D�p��G���c���uJ��aY"W:\�j����(�乔Z��Vj����d|َZ�[n��cD��|��=v�;lq��>o��}��������������yV��IO1�Z����$�"H^���xJ�H�\x�W����ǒL��1j�٧H��ȁe��u�S�KVW�5C��e�,rV�y(�%�� -T�q�j��T�QH��挫�V���*ۀ���*����� �J$�y����[�j�I�з���Ʒf�`�����8��L|�z�sI+����N�� ��/8_����S�Waj�����|�EFP�����>V�[`���1�_H��U$�2:�?���J�����|�w��������>���.���3�$�;6~���ffw��޿lq�����,'	�.,��/����/�_��ֱ�3;�;�c�����?��í��s/�ڿ��;���7� d%�.rl͝��n�=��\�D��sm9�q�"��Z�3�˳ᳮ�7��,��y'aZ��<��̤���o��,Q�V=,9+�$zE^s�s�#=�D�#�	x��}a��a}i�s~v�/�����6N���V��|�����]d� �z��GT���n�w����a����o0���纃��}�{ӬT!{o��a�ryj0�0xZ�A{�̀��Ͼa�	��x�[K�	m���q�v2�����6����ng�c���0H���/��~�O^��y���%�����klg��x�=�/�q���h��KË׾܏��cj:�Q�;.�_��O����?����"�N���׸���fV������`�dƢS}�T<C4>�Ie'��X].��x�e���j����\f��S4*i����q���v�����kΥYX�/^��-..&��7nh����,�̂W�2�-��6݁E�Ԇ3�'�`ȯM��QI1�Wu�9"8���ѥ/1]�*x@�}{)��g6x~���/��`u��ao���k��).�>��LՊz�#�� [d�C�dw�KP����q�����~:�Q�_���%[�Y�BAd {��]��'����1�_��0`�W��%E��+}��W�|R���r�u੕�y30��ByC7��*��'i�,�(X��q{��w�M_�}p�}�G4�إN{��,��py��B�"W�-zL��Gp܃�JL3��K�Ur� ��EU�_X��&|kW�V��8��WY��}3M�#?��Շ�i�R����'vI?�WD����x �_i$�I���5��G<�cn���Vo�Yn�{�Wz5^���$]��4��/�7Q'?��]C�0�d����=|yn�.�F��5���b68S$�T#��s^~ᶕ���n�	!;��]	.}���_+_)�*?�2��el�G�L*	�e�Jy�T�|ބ%[�T����ݜ���5���ܰ{x�s�t�|�z���׻�~����]�[�އ��?���?��ߛY�}������������s���ևE�����a��~�dw�۟�W.��}��d����>��K��Oo��qK���:�驩yl͞�������V��~qs�[G�VOW,��6g8�����7_K?�f���O�����ߜp_��O�9�~6��1���p_�K��f�ݣ���wH����q^	f�[__s4�-0pػu�{쭏S�����%����[w��罾;��#.�t�ڍ�
|�թ}V �sF�X|*�%N��:���܉�
����\���Y�\&ӘY�Uq�[B+���#���p�	����&Q���������D��J�?�����.�.���[/����]1ڋ+��;����/��/w��=O��;Ow��˿�ݸ���_X�~�o�x��?�#��qR2�]�IwL��c r8땤���� ����i-NIJ���ɵm�W'vrv��` �]#��A����}�V�l�;�������#<͙���ai��J�����7 )gqAԿ�ͳ�u��0%q1+<
i����e8����%��X
;I"Jl�a��^��,�N�٣�/��ñ��M1��O"5$MX.��)�R:��t�kx����O^�2�	 �ޢ���Z=��'=kFL#DD�§�Dl�]����L��6a���|%l3��_��Ȣ?mk0�H@���?K�� e����H&+ER��*�J�vL���v=H[�K %i������q6��5�$���i�\e�}��668�_% �׾��؎�D2�_���,f��&?#p)C�&�r5'}�/���r�9� -�[?-���M�/���hE�����xVUg@D���H4��AQ��rN�U!��Y	[��72��ˇ�����$4�������S���L�Jf |h��(�B��X4����j0��	3c���h����� W�I�� */`�����d|Mk�%Op6���
��+�]E��*�6$��Bg)����g��ž��5KF,Pܾy�73���O���޽��Ǻ���w��W�3ݵ���;�o��Эq���?q����\J�z�{����鳗.\�M���}���s�L�l���2h�(�.��/�Q[�1�[��Wm�:"�qQ
�K}�Et|�u���X�E������|��Ɲ�'��-������5���6fenj�q���po��[���\\[VF��y0J�ؼ�{(�Ͽ8{��K~�=����uǼ7��`�7g����e -л������P�u	\�����[�Ȝ�t�
CEv�;:+}=�J2�z2�ew��|(�h�*��%��(��{����'��1����F�����Y���|�7���������}�����71��6
����l�����?1��������C����Ou˼]�.���ݮ��O�����V�!�<�.�����x�	��0[��%+f���.�`iH�ٸA�}���Ȇ׌��[��R��//.�z��ٵ�u�{�|v�����UNnXf�<'�zo�q�K�T������$2���	�L��P+=��V�~<6 ��~�q�rŰ�O%A�Z��/�H�"���_\|W-�x��iҒ	򖳘�cY��@2����D�A��d1o�\�Ac��P^K7�O�J)��	Z\"E��9��a8��jT��TeHA5H�4A$�RԎ��J)E��������hP��V~"�KM>*��c�H�@�	��0"�pfG�d����f�T%\;ޢ��g �*^y��~lŸ���H���ˠHS��?���s�a&Sy���R�[���/8
�[0s���0���[��yK���q�LUya6��(W'%\���n�V��V��69D1'�BGq��[�:�s�N\1������e����40���
+H������X����@ں�^�bz_�T꿈Y�Z���PpxMQ�����-V�u�F�U3(�D�J5�����+cT��6^���+�!���� `d[`��7o-�	TSe�y���p3��p����OI,8�(9��]�*�ƍ����[>�(���F�wwOG�i�xo�{��W��rc�{��J��o�������[yE���j�o�8�x���jX�8f����ol���~�j��^�_�v�--����i�DF�*��';��b=�j�[ͳa�j���c�r[��*�N9���	�&�����е<L�6|�����o�����Пy�;�q��7ׯ�l�=E����[ׯu/�|mk�����b/�[^Yv�.g��лCU[���觩�i�ݼ�F�t*�}:����
S�g�È5F�B)U8�WU0tF(��gm2�+��|�S*(6��Yc��dh����w渚2�.=�P7�=�}���_F��y�Nw���o���Ի�=�lpk�;ݼ�������N�E���=�/?�����6����\�2pmD��/�������+�����1��m6�.�o{�_8
�������
qo���v(d��j-)�q�+�k��/,-f��.�A����w_���l&��y;# 3�b���ٰ��re/>ۀ�"����k��W륚F�d�ڈ�re>����<��hq�R��IQ̋3ϤJa]=��[8`M�z�"��+��`Ld�bUO���7�D% Yͯ�*����n>�	�:j=�N��e
��m$�\�=��R��#���V�J y⛿d	��-�N�n��7^J��kM��fr��~ȡ4S���/<�F�=`�dI��TVɒ_
��b�Tb�P��q f�:ac{��q/�s���Dyu��U��vE6ax�8�>�sET�����.�+�2(ad��ad����:���\����
�H�I	�0 �%s�t��#�M�pi�J�4y1��U\꒘b�iW�����+,�Z�4������2̓  G����"����S�<�j�|���W�W�*�����TK�
��4w�S �C�i:�)�?[�T��>���/�����0l�8�|%"��~��3����ޔ�L�*�Bs��z�
��S�?^q:Z�7����@3���z}x��_�/]\�y������n����r>euh��t�w���[���݃�_qo��dj~8Y�?��g�Q���U�)ou���g�gH��O��%��L���%?�C#̪��Q��b%�~���[:2W��\�}�oy&}uC��o�Ϧ���s�?�?��[S�+���;L{��q�:��\���\5u}��J�W��~�������"!����߬Lu)��	s
�n�8�PHϨF{�≯�t�xe� ��?F�y1���Z��h��z�p��ƍT�$+�B�����|i���)w`�έu'+3����>��/=�]? ��j7�����S��^~�;�f��ŵng�p�M�ˋK*9׭?x�����_�����^�9[6ݯ]�4L����{̾��n�O.��`Zap�.�ʞ4Fc�S���>��Oȣ��߻OF�|�O�Sd�˴���յ�n�#�w�N�lwʣ�+]/�e�0ڱL+}綸ė�֘8B/b/ �7���k݈�-E�q��7Q)'�eUҨV~�菦�ˢ�ЗX��ZL�h��m�ca Vu�P��c���R R��ңiK|)	i�#3�`a<�H����z�Ӵ�۠��y+�Y��YD�P���1J^��1�waS `�k�R�4���������\)����(�����A�B���/��n�6�Tg�a�ɠ�i��=:� ��xa�f��K)�* N0_J"��t�4�p�g�vG���Ht�$Muh��\l�+����Y�\�D����U)���&>���;��J��_��Z\+[�$��\<�Z�R��e�x�~+8\Y��!�s��"�3e+�J%�_T�"gu\����UW�'c�E��+UV�h�)���ݰ4d<�B�����O�11uI�@ƅ��pZJcB��c�ˏ��K(�V��
W�Y;RR"��d3����g�D~L���Ԩ2?)�.�=�Q�o�?d8��LN�`�K�G��;���W��k��nei�����tm�Ǿ�C6
L�^14����#r97{��y��r0��6R�a��2��]���2N\�X��9��{�Ǘ���.q�|�ĵ4ҕ�صx#&�� ��h�8�^����W�3+l�<�|��̓緎�°̅��挢aX�?�.��5�׽r��+,���ns�F�����ΐ�a�S�$Q3�˛����َN�y9�u�@Tb�͞StrQ$��Dk�ٲ��Fb�|�l�Sm%D}؎���2UeMm)6 �k�'��-\}1O�q����=S3ݭ;l\�N�{�qvd3x8�1�qt�'�� �_z�](����˔���J�5{�^b?���w�-u���ls�9Ž���v��6�{�	��w�!��~dR=�8-FzY���V.ꯧ�0�i��_c-f�*��ƪ(2S>6��:�/���2�/\8?�W���7������X`Ӭq�7���K�'��PR���Fz��(����?�Y8��o|�n�n|�Ӓ�ǀJ�*A�oTAZ�$�[,)��ۮ^�'�z�u؁�X��ɤ��"�����;M.?>��(W3�L��Q�eH�.�t��"��ӐV����fH��*�FY��Ʊa�)?~���o�Q�
�E��o�9���z�t���!���������B'a�1v,
H�:(H��l!��M���+4�?zU����R>-����,?�y�k"_�#Q�	/?,��*M�9� iX���;�k�w%���kYś^�D ���UX�2���H�K_�3Oqr��pi'���k�����*7W�\���fFI�#����_�xSo����GxQ�ʯ�zh�B0:N��;���@T�:t��\�$U/�#���z�ӞD��;�ƛ<U	�5�(~y�
��d�eL��ݤ�d��k��"�1}�J����rt���[��\e�Uu�vmX>�!�V���G�e@U`S��,R	U�M����w叾������"5<��SB�����F왵�=�#�;�c��E���B�Mb�(oq���=б(@���Ġ�r+bk�X9~�=x|�7k�u��tS�<;3�����{��S!qxT�B�[�d�ϓ�k���o���Y��O��y2�ps-�a�g�o����k�ڗ��׏�M�°���,NϬ#PWH�sī/G���۷�m��.i��F3n�� �Tr>�q5BB!�Va�XI��b�
 g�B�ƔFM���Kl�JZ��A4'MM�����W��m�k:F�,h���)�6�ACZ�g���g���ӽ$�U�L7�n��A��*eff��d���xux�=�F+=�y��J�,�pt[�>VrP��YVV��ͭM��������a��s�]7Q�u�� W��Z����h���v��$lU����4k��ϳ��6�c�_��{���veW^?���0g����t�Y�@��(=	��C����օ�Vy�����%�X��=]��+��0z��J+�4|�xZq��E/%`S�U�a��C�`�tN8�3�B?��OA\#��'�\����˙GI����gC�z�k�O&�)|�H˛@!�~��vO�"���E:���R-"��Tb�*��0S�X�L��k�x����N4K�(���H�FJJ����
�[��[D��a�R6E����'m�+@ Gf��Q�Q��x
�Ȅ���;M���,�4JT>���l~�N�<�����df�ݖW���|����*��֩�ɫ�6x����Q~Ւ4�.��
��.	���f��E��oU���U0@�%���#2"�,�DS�h���(���F���T���5��$^j����B�b��]���Ƅg�� Iy��1�Y �	�i����
zm�TP4d����8���Y�Ϣep�v���I( (���7�e)U�MO�\������q��;��+hˋ���M���#2X����R&;}�J�CO��<e��W�NR��+�f2ȄەX�*�� ����E�̢M5O�#�H'�*WK�|utim���J.����-��ҕ���g@��3����x��,m2���?�?syajv�d����������1K��T���"�6�{�ш�:v�Ȼ:3��|���QV�����zl|�<%�B�8K~n���L��n�U�aG�tT>L|S/Xae���T��0n�\<�?फ़3�_��N�Q�vģ�*�o}g�@Pjv��)i�Ϥ���:ި��[���
�^�g����i&5Gs��\$_ ���+���p���F��(�U�}��W�ǽxݰ���3 aF������
�0Yy�՝����Q.� �61<}4Έ��3��v(��q�?��X��c���l�x����E����Ϭ�!D޹9T�W8/
��p{++h�u���e�s]˶��H0��`S��;v�*I�R�]ϖDՄ�J�e�ԧ)�[�Z"\�*�ie�S\Y�l&��-�#?j��oK~�Z�!,b��FlL?Uј)�i��"��[�4��	�S��l�QA�c�|��5w%�TY��D�A,c����?I�q>��t���Rr�����Y�奸�e�~�n+"�:�
��?'_��a�;[6�33w�b{t�Y�=�wj�5(��$(4E��'屮��n۷!�OQwEh�lW�)[X �yąK��&�Ĺ�������C\	[�fþ�M,d�pz���l�$���}�-J��0��(�=�D�B7���SxO��C� Æ����E�L	P0��]�&5~����+�d�J%"�����	Ŵ#�u��%%9�#�+����TG������O�W5���p2�P�.J(�W�������Q��=\��w��]����U��
����h��&��hIء�:X�d\,���k�J�l�eK�-0�"�*|[kZS-�і�m�AZ��y��9Hy�Ƙ�~�}
�������3��#�4_���|Pe�D�0�������a9i༥ni~�_���4�~����G1���Gϟ��c��d���&���Z�*�o�o7�s2��-_y���9ӟ��w���}�k������s�o�����s�l�����Y"�~�+,��qm8���O�_�.���6�s��y���n�e(��Y���� *�k	b�N8�aa��ԁ�iY&�D�|
�-2T��
h�QS�(�����
��r2�1�=��洍�fe�ʂ��f��sx� +�|b�m{{���D懩#�,?zH��4G���~U�������[VҎ�^�<��������U���D\I�u)W [l�s�q1�A3�Ӕ0�0�þqd AC���i�}ee%^=���k�@�Y0r��\d��[x���2��̹XEn�bXB��do�^>i���;���s�Sw�Y^���vW�≩S�tw��ɗ�OM�c&�|S��/�lL)����bt�y�:u�ơ���|Z���q"��Y��G(S�	J�$����ԃ�&��&Oh����$U
��0^�!�uYi$/���UH_m�׎��B 4�6���B���m�̖/|?���%?f/R��;��#DC�a�A
�w�l.�؏��3`��,S�s�?��~s�3���q�V�������sĭl�^�3��D.�N�@{�e�m��C%u%9��ݛ��->8K�!�x�}@G g��F�se<�K�}N��)3�@�����T��3�PW��R�������Nxu V���K�@��@���!���+9g������]�s�/�%�c�]y�^($�+�e�t^Gශ8Q��2�Y��<����_u��y�ϒ�S�+<��_�I~q��҄+Ĉ�Nx]��$�s�(+�gU�z�B7<xV|�ˏ��Aӕj�v��jس{#��3��R'�wL_\��Q�CIQ�Z\Ϋ#&}��&/�	�O��G�\��?�H���8�b�o�g�a�M��"2�C��l�љ����zv����d}u$/��+.
��˂�$�߁��/o,X%� �}�^�{�`�精T�:�&v� 3]��9�/t
��o0�#�Vl��ڋSHI��<&�p�K������������������������7��Gs����W�o~�o����a�(�_��8ӄ��e��������w6l���?�ą�����e�������_=|����;\KKF<��͢+t^lB���@��[.�����|v��5���v���CM��r�[4��\\]��:e��e��W�-�T��Bp����ֈ��nD����9QKڵ��5��X�E�W(�&�@�vi%g$�e��U?���j:>X�eڹ�m�c�LA\Q�*b���¨٭�%K#�v ��k:- ��~ci<�q��R��(7�����a��)F�W���FvD���p�s#?�zL��o�:0�(���|}�---��%�c��yڤe��hXx��:+ɰ-W����<&����)�����*�,�c���#��3#!3Ȉ/^���#bP�1��%��8�P�����,�-�<���`��?oU�M3��r�s�O���Z=M�NB�v�v�ff-"�KA\aa��h+����F�2a�b�)L@��G�3Ҁzد�QP��ZE��8Ù#SK
t�.�G%�f�:��N�E�5�9����N�	��%lE@�i���Í  ZIDAT(�"��'�/!Q�5�[i��0��u�-��s:.E`v:�s�����oߏ8q}}}v��aq10���0�?�@��i:w���`��1vD�a�Lv3ؠ �]��:Y݆�p���Nu~�b��8����P�9�~� ^�@�����d�[ ػ!.y�yC?B_X�);Gat\����gꞱ�A��:';;�`s�<Rl{9�L9h]^X8n�����G	��Q��D����y�SW��'Y'�G��^�"��$ݬ4
砚�}���!U_x���Jӑ } �G����z(��������}�u떼e ����R~�+y)�e�>Lw@�ߝ;w�ĘA%'uú�^t���oWm8��v��n��-G�d�=�x�A=@�p�Y|q}���e@�vk�u>�˺o���;X�kl���o�ȁ����;�킃$�'��U�b�K�F�����,��oX� /_�Oq��,揺E�d�(L21�Q8�2��O�����J�HSр�r��񘦼X��@�˺�����w+�^[_Y�v6�'/?r����G�v���W�>��X4h���d��g14\-��_/͸�t�7�g�ټߊ���P����a    IEND�B`�PK   W�dW�Q��� y� /   images/7a682d23-8f26-4a7d-8a92-f03913074d3f.png�{<S�ǧ�rY*���B�r)Y�6׭!�%�>�\+��!r�!��2��_��ܦZ����bi�n����s�s�s����z?_{���Y]?tP�   8t����� � ��!��jww�s�% p�  l��� B4 ��; �^.  @j���{B�.��)`����e�vG�߰4����t\��+�;$�de+4\Fܝ	p���m�7��_��ΐIL<���J�����]�>\��F�y�E�zYQ��͇�;�����u���x�`
rUܸ
i}@�7�۲�_���h)`R��b?PY�vMm��'U���;VQ���SK<���g�͉�=q�T_��A&j)�c	�X��°i��HR�}�֌�V�K�1`E;u�C�%C�.�*4Ǡ>eIm�Ž�fm-R�����hX>��:9 ��_}�݅ ��v��5��_;u,�A��S�.�[?�8h�U���h{L-s�)�ױy?��OR���0���\oS���R0N0d-���+m
>�Ci�S4/�D�N�l6
�m��qK)��IM��n�_��� �*]�CZy��<���� *K���S�P����S��(�Ts�'p-�麀ڸ�c@��֟�f���pͧ��ERF�LX�=]C+�����b�ش���P��1��J���Q�dQ3��JNZ�	��VWC�=�}
B襙�B���n���F�&�Ȍ����	�%ze��Jyiߧ{C�GT���i��zE�閒�~l���{?���^m��
���e !�7��qy���Dˬo��3�lP
T� h���}���$>�Cg���~�X�
�hb�ծ9�2C|�g8�u&�"T�v�@�_���o�#H8`�hoK�8�+;��YC̮∭DR.�hL��@μׅeլ�#�������@'V�2��'=��h�(���[$�t�LB���fh���4������������*�(��:ψwk��������0��/��5��b7՞{BI>�:@���I�J�:Z�!eͦ���&�9����W#y

�>��K�#m��	�t�2Ǣ��:���#v�d��w�ھ�Ǵ-_Pi��'�T{t&� ��Q�p��:�T|�tȺ� g܉*�c�ޱ��]:���ۜ_�?��=��7&@s��!m�З�1??�3����M�,�^��2�*"{A�e��_�+�^��!{A����J�1M{�t�;9�(kιw��kf�ٻF_������BZ/��1����J-�J43�8u.�1���v٢��f� �ʫ�G���5�f�<�K�Sws*&�}�2�� ��^ �R1�)#�Tŕ3V,�Z�C����B(��^ڝ�K�&�@�*	�����R�ld��|�+8R<�ˢ��La���ZNê4�f���Q�Ǻ2F9�M�������/�ʯ�m�����on/.BK��t]SS�ֵ�uڴ��6~M����%�ſexht'��T��]g>陜5 ���d5������ =L*Mg�MyՏN��p++A/�|��$ ���A0+]n�w�ի�B�������գ��2y��^ߚ�'fHmՑѸ�C���T{A{��؄�9�-VeZ~~���Y�֏��^r�F�'�;�,,)�W<�l�������A�8­ O*�?+�s8��9>N.~������v��>	�:$��[DO�[¿(�d'���,��@h_aC�9�`'�>.^�'KQj���i�tUH���Ҷw�z:\`�`�z��dJ����A襵�������9K��!���!��z�OȬb����HI��~���l��Np]��8�-�q�d��a������z�Իd��5��qƌ���(QK���^DUՕ(�mc�L��n랇�`��fnM씩/kc�ե_č-�}��4�V/g�  Jk��R�n8��~O��v�e��U�`��ê��xp�[?'Ve�q��+c���i1ˣ�0��
�ubp[C{ހu���ܼkx��qo�}fA/TݓN�<�����F�Bh��	b(O
�_���8/Y�08���}X�/H�ZP�]�=����=�2����'ͧմ�(q5P�4 �	�<��`\������S���?|e�5���W���ז��T�_���W�S�~8:ߪ�Yώ�Y�?�
4čSK_~�~d�d�9�	V<���׺�ѷj��ѕ�+>��
���	K��.(_뉢���{D������w`¾K� �^=x��98�X�~9��ك�c�J����(���,�F0������EX�Ad��z����JE&^*�?[�v܌Y0p�4����T73A��P<�[���ϰ�}Ƶ a#�>kg3�;t9�6?�g�L���;oP��޾��n���9p:�ٍN�?$,��tF�щ�J�9��ia�����*����I+���ĘK��p� Z ���Ϩ�L��xR�уL,>���S�� �|:H8�\�[���ǟ E�~ j�3�y�FX(׋��Q�*� T���DAs5c��'Ȇk�mى��&Ý�'.��.�e�Q9g���L������v��B,��p+�o��6L$�L.M7��z��P��{���r�zz:�ڳZr�.R5�V|��)ڮ��@b��:z���EhI�jj	?���\���y%��y���~�:�ϔ�C���E�U���lR��砟 ���&��R��s��Y-R�p�q��RG�C1�V����P���FZe���+)���h8���r�Ӡ㏥��Z�P�����t�y�S x�i?~q�V�,�p&\���#�� �Acfz���G�-R偖���{�m�Z�+�����c�X��%(��i�0cf^jsr�j��< ��k�[4 u�A�rr�d�;su}��][y=��m4q�Yp�g���zK-�(1tHww�5�RDb�3�	�?>�(��`���1� �{pHfVBiн����)L�Ok��&��G}��������+ֳ�{�FoS$���q��?���ݝV��pU�
<!w�6���\+�UO����n�=�)1_�,Q~li�1`^�0�S �bn��쥘�G��A���dNġk/(M�X���+�0�׆���[�D{��*{r��%4���T||�ώ�R�t�}�����8�^>�+ª���s�=ow�5T�V;��ب+���z
<pq/�H�?Z�w[��O'�=�u0�֠[J�A��OV6'����t�bW+e .�"���쉫�co�*G�� �>�� �0��{+{7��rVv��xa�����#�R�b1��;�\��t1̗s�d��%f<l����q&8�i�R�hQ|XG����2]�� �! G�
屔������������?�91�A9��	�f�u^G��nu���!|�&@�#����i�uN_�>:�h�����f3D�D��L(Z�}Npu��8�;�A+� G{�G�#�[q��������^��zbO�G.u�6_g�U�/AP�FwT��uS�ݥ�1�X�/��~Q��~�0!��Z�پܵx�y�7V��ɣ8|��5���p��+����)��Y�^�m:s}�$�*RU=՞'wZ���!�~�2K2����"��ڸ�M�����B��]x53�:��\֯���z��;��j2�����NH�<�O�9V��y{	}�Kf��M��z$�Y��А�yIʿ�Gt��Ѧ����Rp�r6Ho�cn��I��
ך:~=Z�m�!P�T�t�ѧ@V�_Ug'�w����G��q{�(�K�QiZg�z·�&tB��a�M���q��Gk_�=˩���3���eθ2^���TB�V
p�'Ӟ4��]��kK�D/>�(^,��� *�x�yG&���tܯ�-
�����k=f��Za����R[,u�b��.���+�B�m�2>��Pz��R��6P?���v�@�?�t9�4㱾��]V|/�~����h�:���6t@$�Y�����
W�ф[;4�&��ДGW�����)�S�Sٵ:����6�6���pP*������7�c�/�^�p}� �?2oG�z��ν�\2�K�e�1E^�C�>�(q@�u�������������^n��?vg����	~/�qW~�}L����գ�m>ݼ���3�/���킛ҟAϼ���J��r?6��[G�x��j�����^12����Z�����UK�Vo)��kQ$6�&�ü���r��åB��\�n�y�y�"�G�f�or��z�e�/��������b)q	���v~{eun.9��K���Ⱥ�mm��j���f~-z�>��z�O*{��o.�d7,���V�c,��W����n,�٪^ ��������%&-w�=T��,)�e�V������^YrUԈjo��J��&��>B��X�k��-�t+�u�f��þ9A�e���1����}8�T��κ��W��VY���f�����O��n)�a>�ѡ�KqN*����T�荑}�`41�S�x��`�����u=~|
/�9!X��X�vm����Z���ʔg����En�����w�Bg[�څ�Y����m_6�<��d��;���g�Ǆ��)5�(=�]��[I9��7aG�/w�7����u��,�z6�h���zj�����φN���-��	vrq��i8�v?�3d6���QԘv��WXJm��t����c��E=��u~G`���k����p��_�[���xM3��F1CFa'��.vE������+���f�ؗ����N��3t��������j�ԶM��)	�����>�zp%�z�%C�Ł&@�����g �[�]���3A&��V���h,մ��f�xh�+��g�>q���C�Q�D��<C�[Ϯ�����m��ݶ+�8�&�nz�<��jDG�B@S�?%C�{��G�`�����:B �,�\��;Ћ���@I����� I�"��{�_���Pptb{y��R������W��1Y���̮�Α�3$L��W�ʜ%�V�tݗ0����k��̳���.�]��3/x��0Í���K.����s.֗#I�N�W�n�L-n���ߎ��j�����}�#���I��O�?�n�3�ϰd�ŵ͟�|o��pK��ti�Lيz������މ��ة�X�l�B�z�J�S'��n�>�hn� igRaGtgq���C�i�!�i����U��A�Q��pRC�g���b6�)�����%����.�8�l�N�ٶ������J���D*�ز�IP'��?zYok�p�s{�p;���T�zh�j=�7����b��vU����쁺eA�����^�E��'��/��p�{ɓi�d��@R��/V1#to���ڊIP:-����Յ�cLb���%�+��j�F�˿ (�A�<�ٻ�Hn��C��.�-�F��X�v*��YU������n}`�(%���3?O�n� �_I��}l������_)`0�5�W���?kSl!�4�f[!�� P��Tiι�Ԍr�����I@q��K���'�E��++Ƕuꔸ�w�i�G��n��ܠ(D����b������)@����Zf2�s�2�s����!ʾ����5���M�ʡM����ֽ�����x���t~�"���Η�m��q�+����q��L/�}ҍ����e��r,胃�Z�'k��7�fW��eee�?�+�6��8���p�����_Q���w�h��@Є��"nĲ!�B�*{bc=�ߵQ��Y$?��-[\ḨO�B�ٛ1t�:�N7���2��Ϛ��Ų�&v1���磓q��q��S�0�%�cs`q�g�/$�HFq=���-�˦(���}g>]E�݌[m
��B��4�H���� 9�o�6�_�u�Ǌ��3���w~�l�'A�l$|=�a�@���XM)���!nk!�ٚ6f]�K$c�P��$$x">����$f�d!�Pp:-��E���Ykj����g�1�l�4��&��v���5@�xk5��b�k�{���|� ��#1F���'��<� d�(5��(~q�#&#�\�YO���z���u��I��%�q�}�wpY��
ܙk&�0]B��a�*6/W�������hLߐ���8L]���Q����VA���yt��lS����&Zn�|�����GzZg���s�Y�n�)�ç�|/�N�aQ��m;Ck�k�]ܵ�w�z\:w�@e⩤�_ۡ*!��0��+��g;�|�Ο"�g���4�5�b7R.��x���)�;�H��+IGG�Z��:`�����R4����Gb��s�<Z��8�����A�Ư�4��{e����J�\�I9ܮZY�����\=�nC� ��#������5[�zV��0^��Nl�ښ`�Tvֻ�G��v�'j�t�UPIG�-2p�" |B��S��EE�7��4k�s>�/z?(?n�┗VBp�G#X0_�O��W�}�7Eٳ���ۏ-�zί��g?��H�[�G��27�ׅ�C�v�T'��#iG�`�1��58K�Y��߮���ީ[G�7rS��:��z��q�0ԣ������o�L��>���K� �/k�䂝v~JH�Y�+��S:b�14��X�'��Z`{˷�k�Ʌ�t/Y�]k��a�'�FA�y�
���c��g8ݰj��)W�� }u�z/vʋա|k�j����G���6��8l�dQ��*qWE�1�T6�;?x[��[l6{lջm숀ƿ&�����1.�_�k�A��n���.c����Ob&6�K�-����ڵ)���Gy�|6�m^�~�o�U�O�]��ĐJKz�K$�~h�-���n�`��{97����=��NZ�4�x�-��k��Q=�;"�<�:4?�u�_�E�l�Q6��b��u��9]����7�W����lZ���)�d����³2����|�(l<D����VS-��?�ޝ[�^���U���VU����y���7�b�>��C��T�lJ��K|��o�Xv�L�5Aii�Q�8��f���TU��r�6�|�O�b{e;5����p�o@ty&@:r>�2P�m���X9��e�� jK���I^y����P�C���]:���m���8�/Ŏ�J�������k�g@rS�r+�I�ʩ��)�ϽK���F"�#�뭑���
c�C�Y�O��撽f[�`��.E*|�uk��;�ֶXQ��3_��&^�V:Y,���YY�c���.Nn��qJ���{}� ����Dx�ɀܲr��Z�k����u;�Kg�KgHf'��Q�͛�����:S�)�F��	^�{5x�}�׻Q��y�?S�ڋ�/s��|������Wa�ǈ)�R8���,y�T���?v���~�ᴤGa�^D�B�ۂ��Ą���A"��-�ҰaS.>���������j/bY�
O�іWV�b)c�N��G��!ͣҖ﫱E�]���y-�G%��U^�Q:'�������%�ИG������߿{���
��0�x��j�r���˳���l�ni�t�[����������\�qj�L>-	b%����g1��r[�{F�����F.�ss�y&�^
T�3�RKN����;h�#�x�}�d����/a��������hc�i���5�s�ac0��]�n�Ʋ�^��WN�f�^��f���G���}ڴ��d���8�?�T����k��6�9q��o�ͶOF7���5ׂ��ur"��)�D��NU:�4����mai������>�S9%KMm�kk����$��:&W��Z��O�0��o�6��lm�� ��b�@��g�t�dk�3Aώ�M}^5!v�4���AU���������^*"0lϳ�n�{4^�6k ��Ռ�+�I�emX���/�h�����E�Q]���:�*P�R*�����>-j������ÿ�;��� �+8�:��j6z�7\_�u���$��;����5!;�[�}N��߃�_"�p�#�kx�w�6���
����(�FT�*��8��zg�A����E`jEyy&�ſ=D���jd4�;����_�W��"��@㸱�S�-�u�W�Y���
�?l���zW��u���kg�c�pH��	��TW���g��L�\>��/�'��9�:������[���u�­��U_��I��y��K럮+���:%����:��R��ʯ�%Y?��]j�H6@W��F/�D,�Ոy�X�g�-��bZo`0=L�K�V�2�,rÛ�� ��X�iB�r�Y��X۰a,>P���cY7"��~7m���l�<^���?��lՆE��;w����0���"�!-&��D�`��t�˕R��+��k���S"\:�\�+�On�GϬL��b;��}���jZ�z�K����Gol�N���%���.����=&��s���'�-��<���12��<^X?��ک�z_P�m�3�)�T�na�?S2m��7��))Nm!��������?T��?w.y9���M����.~r=�Q�ۂYÝ�2/L �?�s��l9u����� ���/;���)P��T����r��K�<��'�fA��M���$�^�n������Y�Zj���<���fV�R�Q"厖nͽ���=y�'a&�;�'��c��nꞐ��r������ԏ��h�n��L]��T��ǚ�K���t�o)�DT�L�n���>��(�&��i�'��/��mL�{��� (Z��N�3*-�Oe��-E wn`=f�mONֳo��m��G�����um�����]�A��f�&g[�}�
c�9�c�!�)����xp���L*�=1J����[�z�噽����1j�={���}q�om�)ţ\ؑ�Ys������K�t�?����r�N��ƒݏـ`_�����J_r�rAK�^��~zu�(��z��>�Ę��w�����IIq����jőK�*��.�� ���fw��?�������9�}D��G�C~���jx��C��`�9�;35;s1M������E��).�f��Z,�d��~��� 6|ω�R�E�����	t��� �V)'US���+KzI��/�!߉��G}Wc�- �{�ү����+�6N|]����ċ�E�>O�W����ΰ��X�o�ڙJ3�\��^|�Ե�5�"�*��� o�򬖳�V�R��D�S%3k-UK�aNK��!.Q��~��(���)a��32���\Q��C[�{6c���ES2p��ghc}�M�vЍ�,��x��mt�*�f3�w��M_���@.1�o+¶˘�{�ʿ��q%]�L둬T0��dճ���{mݳ�M�9��n3�fU�&�<�(VK-�)V�bx"fe�]�s�qF�C��:�3j�h�k����n�6��5�W6�Zyzo���@������`b�R�u�q�a���^.�*Xz������[���_�n^�((�,����
�+��[[��^$�wjrsnd6� ��sl]�D�R��=��P�jn-$|�2�6�?$�}�<е�/(��y���o�M��9\��QD;�n>- jNC��%L�p�� Wo9��� ��~	����:�4(x�=�t�<r�6�EjZ&�mv� h���d�8������=wIZL�.��<��7���ekx{�B�����J�t�z���?K�Y��x�����	��Z?>Q�vd�/�Af������e_�n�yҫJ5�N�%"t���M���q2�ރ��>�8E6��C{�����Df�B됇&�W����_�?m��W�����39�<�l�7m�Ӛbc^΍�cE8Id���D�l$�J����0K�r����EF��.]��\z6�ߍ�J�	�F��M@+�����)u���Q��bo0�)��O���b`&���9A$�н�a����s��oǬ���,�ޝnd8�F�
R��>�"gegnx-z) �DoH��'�&+�g�㑚����P+^����ƚߚ3/)tDܿ/�h�A���x�cT�x�i��u��s��/��@/0Jnn���Ȳ�����~��
���N.���`ld���R~U�Wp��"d��z��3��t�k�PHH®��ƅŲ�N>�$u�M�l��v�wֳ{��*��{ތ �����m-D K��� ǈ�����٥^D>?��=Ol�l)��;�P�f��[�U*�᲌�C���e�ؤ!$������gX��3�������4�����u������%�M���\�h���k�� ��}�ʓi'du���:��S�����n'����P�O�Y��1�z�ʾZ�����I[�^�S�����]��"�	����D0>u�%P�8����V��D�N�9��%v2�,j3}f���<q_�/ķ�~!����a�XU��A>y�pd|>�ԧ�ލ/yנ�t�:0�q]5�OtE�D�=��iw��S�A�DKX�+;��:;���a�(-��c9�q�eRщX�д�Δ[(�����zm��5��io��D����G�����ނ4��f���/8E;6�Tu|�DQ�A�����?���w�H��9����W���V=�Zd��:י(�+*J}WaGѣd:���Yp���{r:��n��!�d�sӃW��B{��p�IX�nraJa�M}�83�g�kˁno ��d`�j�t�����8�á3���ڪ�������Z�bg��9�@�X
���d��N	��mf��V'mI�\=}�$��p��_��ȏ�3�υgܑ�C��p�>�Gde{{!ܑ�gS��9㦨g|$�K���,��{��;w- �k�Px�%;b��{�=�s�dZ��CZ׹��B�x�U�w㩰���<����z)����.Ga�t�y,��'�!�E���yg%��Y1���'d�7#���X�xs&�d���*iř�C�L�[�ЪLe��-s�Y�$�n�rP�t�Y�}�΢܋���7,��fS���Ni�qL{���n���J��T�D�X#�qX1�6��^=������~趨�/-���~��M��O��䗶ee�iv) a1Ў'�2�����2�O�ϙT��/���2�wR�}�)'�;z\�i@�A�W��Ua>��=�n`f��D3q�L�����	�URo��j[A����
�=45\�8�	K0�34З��@����d���7O`����%�vYS�S�ҏA� 7Z�KG�*ȉ���3����n�	�w��7bGzmء�_����Ko��׍�r���{N�<�����B��Tc���>i��� �666���G\1׻�o���E�h���/܄8��D�_�h HVe1�9������M��=���EVe4���_a�}y��� iΥk���2V8�D����H�8&�؋���ːv�-_л?]%v��T8�n³�h��Ok'��¥�h���"U��kb�r���tHeY��|��h���W�������*?���N���>w���o�NCE�5%��zx���Us�ikw��n�=�����g98|c�o��'ԏ��a�k��ѳ�Zx'R��Ld���:�h]v��u���͌L�>��1���Kl� ��_��&
k��� =s
�zv��>ӟq{o��;	L���7[�z�:f��Й��azY:J�'�U9��=�@iq i�\T>p<�*ҏ��j����bu��C)��-��h5{%u�\�fN��T�/�7����$ˈ�$��j���`�bgJ��׹�������\8#�soN7�Yi�����_�벃����idRif����N��x��|b��&�:��CT��.�ӑG��� �2Dr�=!�X��ӹ�MC��ڨ�g���W��~��BЎ/S��*�����B��G�?���~_��X�7���ξ+QP?p��_~�W4P]xm!�RQ����#�g`��qyZ
�{��}]m�m�:��C�ͪkj��,ـ7u���E����@����$q4%J�H��72{v7���������L)I�W�!���ʬu�c�P�sT�������ʒdX��dۯ����B=ԃ���Ǻ�˧�ąt���R����"�U���[ڹ���K��y�^"��	�F�����@�7@|��@���Ĩΰ�Z �V��ţ��{�[2N��~M��{�:����x��!�X��Rf"�����.bY�^a�#����;��98}h�ʲ
�տ�66�q��^]��BH߄�*y�_��ndͩF�}c{���7��͏9!��g�
��ǣ����V�K`C۴h:<x�4���jda0��a�җs�6�l&�����'�z��N���"�rw���q�w�QsƊ��-���M�,|��DG�7��Lm��Eʧ��%���B�U��J�rn�|������e[�K��� I�ܷ3K��/93��`�,��O������q[Ɍ�g�)��Z�Ύ�l5H5�l���rN��=�Eg���f9�6/yJ�xd�4�V�C]��m�����#i��:�ꐭ,)�<>U3��$<1/��Ӗ����t��h�NA��q��<QY�O�}�0�;tp��f�>�Ǚ�{�6J�'�4�
*���{��/�vO�oU�꥿c�z��{���A�r`;G�ч�T�1`�r�t=�M���r�{��cF|����<[�f��b�oNi�p��_j�RCr��vW����>1�B]h,w�5*m<�i�${͸+�7}%@K|b�
��[uS�n�uÜG���h�]��:����S4����k�Uݐ�#�V*��J��q1^6�}��__��ɱ;�M
�f�l�Y!ٔ�!Uʜ��������t�"��d�$?����f����O��t�s��qՈ#I&�b �+ɭ��E��O����r��| 	?���v]�����H#E��K��JH�'�@e"H]7K��W�x�to�fz�-	(^y:J��&���q �S� ���Y�F��;'m_=�RV��ї_]cgUfCٍ��cma���ҖG�Re0yRYzetk����o�U�ږ{��Qh�k�5�9W�\>��<w.���=޷�����+O����^��M�&V=ɁC.L��n��y�_|iXk�ȋ*7yZ�A�ؽ�Y��w��O:)�,-_L���ZWe#ş�ܵ!��Zg�K�d~�򥄨��͞�g�mS���^$ېNu���D�u,�zI��%��|ZW��'G*���.Ą�|(�m����h	��eQL�*���/���6U,��FB\�嶢8�]1j�d�Y����s�n��.a����}�͆�Z�p���#[���7�F�!�<Ӝ�'�A=���N4�T�BΘ���p�2�^"> �H��͟�"��7�-���Wd��!<�f)
��M�Vs�M�!��1���+W������^���������v���U�1� ���o����VF�uw�-����N����	��#%��@���U�������%��!�9w�{�g���=?�-��˚n2y�F��"��9A��LO�Uu�"�{��%�h F#��Vǚ���j�;�Y �ͶX/����r~D��[W��u�I=G@a�w���)�,�I����k+��Տ���1a�v7v�Us���2�ԗ��z>}W-����,�?�^�n��DDx����8���ea<�)�w�ۣ����ؗ�D|�Pu�D�ݬB�[��Y��4���Ն��+;bq��_��X�4��2`��%D�  �K5��r�~J�,���0:����j̖��6F��A	i�\^13�s���Q��{�@�]7���
y./�ca1�?L�����"�ܔ��&�]��P:�|d���z<N�Q\Cg��?�_W��ŖUW��(�|��7 zU�&u
�k\�ef�v\�R��w�:��"����ug3�6�U�cu�S�=��`��܍ Nk�II�	N�}ܿ�I*�?��!u��9�N�4F�����7�i��Q�Oy�sú�?xtaN-�q@�SB`���CwD���W_R��x�ΟZ|5����[N�俤hӾ62�:$�גY7�������+/�����&�	S�L�-�̿��{�82������Z��~R5։��Œ�.����sA�*�Gk5����"�L���[����2��/��ԫ�?�[z&��o��v��LAO|_����wZ�ӱ���~0��"�w$�3�K!ՀZ2{[[+�����U����ªf�=#s�!XJU�Ky;�>�3����1;��y�7�w�� L|W~�_AS��s��~[HD۫�x_�ȟ���8jQG�ǣ~ԯ)��8���2�X�<��a�=��Ğ���ntr�����qV�_�������W&;#�[����tȨ�q��}t0k�֭ǜ�*�^Z��l�Aְ*���5�o���
)u3U��R�+��9�B����8X qG$��\Z(E�G�^�:>�+.aAa�.,�}��䠸�1z�˕��	�U �MZܮK���{���(9�V_.�J�q��?k$ط�c�])���3,s�̴٭i�����}���*k�k����Ze��ֿ�����+��PW�x��Y�U3Q3%k%�7ʟR������4��	��b[jg��4Ƥ�E6N���1;7����o&4�ѹ97��#1?Я���<�B�}�\5���x?��P`{�����2�)?c4C~PO(�'X�*Z2�7���`�����/��� N7!��� fic�K��5M�M�*�DuI]{�*�:c\Y��i��a��R��/!�|�G���	��"p��OU���~�̸ex1�Ov��~�����ZH�H�bJAzI-�����D�!M���f�(�	�����w���o�>Խ����U�IAn� E�7�"�\+�F0O;���#ZBE�=�ϩ�F8��߿��U�w��j�O��֏gO������@�VTb~�1�eH����{�UzB�m������Զd4B"�c��������s�_�;��~k�ҥ՝X��?UX�ȡ/%ˠ�W@�0A�;9-H�}�o��Vv뫭�������C��o7�^KE;����Y�V/��tR�(��7aqW�|��HX��@BAHr:E��|kr=i�aC��⬓���>�qmc&�K��AY�/��l��yU�#dE�o�S.��X Mjb�Q�/&���Gv;Rר!�Q'#Q@��]̎�V�dhA�ߛ;��:^J���}�����G�-&��r������+��F�J�uYb�)�Ǣ��ɪq�>�X��k��U�4���|�B�J�����ҡx	u7z�@K� ���OC�NJT(�g$7gf>�
;������f�0h�l*�D�b��O~�[I�be8�%jÌ^ʻ����C)8L���G���XR�C��,�^N��y�d�٠���mm|��@��̒� �uE��|C��f��ʢ g7Q;_,A%��W�����+Tº&���rs�9Z�H���O��d��T�奲�����Grf�5\b���RA=��4�Z��A�^�7����(�
�RJl<�|�,�ӫ	������������#+�l��E�$yN;Ջ��5B,ըt��T�@���M���n@"�˼�^ܧ�|3��F���1�u�t$/���KNm�i@�,ׇR���{�G����y��*jh�.��e�Y�Z�=��@	���§[[b�,��;��Ǐ��3ϊ8hQ|!q���X��<,5�ܔ�8 ��H�kmd��	��eyNf��.^��	m�-8|��W����^~�w�g������'�ga��)w�\A4%K�NȏPN�����>w�-Iɒ�W�5���;�U�5���x5�����?�6��9u�ҕ�[���@�D��U,_nά�u!���<����[F=S׳oթfA��Dܝ������wih��#��iq��O���\Ţdadz���mvʧ���u�X�%h�	�C��!��Hx�t�G�'��%�����3r͏H��.��Z�C.�y��Ess�RV�O�����k[�M8��랮��}�����~Q�(ejU`�hGRO�����q
B����Zj�v���g�� �ʼh�	�mzc��_��,ګ�K���GP����Q7����z���1?�w
hTj�9�c�$�/%��Kb.w����H��J���*�Ԯ��b����'bN��hyw7�T_�d�/���1��e6Qq�f��)uފb����������oJ�%�[78��V��dO�l�=c�������\�*=��t	^��=�\�_����h'�L�YlO��}�͹�"�����k�	�̽��5�釻�I�~+O�9���d� ���B����S9����V}�5��|�:��ID�'���zwz34W�`��~�34������
o�g����
7'B	,�����ޔ���x*uJ��w<[�ǣ-m)*T�*Q+V�l�Q{�Jl�%6Aժ=b��E��"�(j�E��D�R�~�����罯{���?�>�<Iuȯ�n'��Y�	�/��w�E�siF��}}{��܆:d�b���+��pc�B���9�w9<`]�S�]
fm<�	̒�?;<�,ٔf3)��],W{g��'u�O��x�s����/�����7ݯ��Z�qn��o nq�?����녏��u��3�R>:�f�1�4f�[�5p.p1P������J28��J�^��Z��:N��W��Ȩ�O^	��*��qmcR��}a�~ooc�/�Vxj���f�Z>���_e�[^Hӫ06\ˠ�q�	�u��4�\�p���ʿG��Q����a���
T�������<,��SP��<}���x/Y���������6'kq��wn�*�N�@�e�A��T���_`3��{��sʷ�d��i r#��ګ�?��܈�ҽJQp�4 HeX��)׭I�Q)�,W���7��C9�L�Y5Yaa�,��ɬЈ�kM�6���Ϻ�Lo}̱��>}�m9�d�1!�tԷ�Ŷ�+k�e���kKf2\RDI#E�Њ+����α����CB���������f�2�1SBl���YZ������x�6���.S(�<n�V���y�>z��AI�K"�%�n��D��(ם?��Y2�ƃe����'����Q>+eȫ��;�]iL����1��rR��W�m���YB�ev;'��H��E���`�_6����,Kca���R��:T��+y,.	F:�z|E��6�P��+��#K
��k+p�=��ɐa+ӳ�L<�22af�n��<�^�y߷�p��,l��OX�q��Hͼ�#գUr�/�+��9�^e�N�p��k��)�XY�$$��G,�兮�өos�0仢I?bP�PK��SM.(U٤�:O`��u����^�-�v�w��օ�!�ۘ�]a#�h��0ݲ�0y�����ۮ��Ǐ�w]���=�X׷^�eqr����M�=�q�[cOti��sRz�2O�+c�8�\���
��ε�����Q.��q���V?�}���JO}�����l���Y(G?�ݳd�i�+:�
!j�]�p&�!��P��K/�ksn���gɈ�{����ⶈ��%4���Ή3��7�IB*B�3���T�����53ˍ�}�)�[X�����|���_��c�/ƙ�ft-���]'-����t���8𵩑�D����ύA��g����̹�������
�o�}_w:�7vJ=��OduK�G��T���@�mzqhR��G)�Y�\w��T!�79cf�41�)�ϫ�o��0��=�"Q�������76��|�k���G֔�"Ȩ]KZ�Yz�|�,0����q�\8�I(C_�%�_~PG�(�E ǣu���<ڤ=V8��s�o�E�s2�f�����-�G.�ހ��C'�3u;j���j�ʑ ���(Hd�^^�`,����L�[���u��޿"�Yc�o��uΖ%�}&m�d�(m�Oz�tƈޕ�D��j4�)�[k�R,1�[ �Im�%���[E]0�^!��W{~��K�saaazdMŕ��?��gx�� ~_�{��T�.��>��2��.��F��i��`t
"譹�w��X�̨gyk�Q���4�,���Li ���m��T�� ؿ^֭��+��Ԁ⿜b�-v��?��x"�Ύt!ydk�AJ�����]�*pX����>+��0�t�y�i����E�X�"� ������Q�F+���۝��2X�{p	�*Q��̓�<ܗ}kw�N��>Åd9�M�Y[�r?)4ό�!�7������a�לh_��g��I���T��F^���)���z�2�fwr��S� �fT1�o$`��/6nf��]�^��N�u��R ��R��73-�q����4�dY���wÞŖ5(��ń��XԞ��-)y�ߍݕ�
����������ں�GFw���.�X6Kv�L��d.�,�4�Ek�o�<z7L�vT��!��n�[��s��X.O�f��<�N|L )��t�����ߏq�*�ՆX�:c3m��Lߎ���D���4่�H5�I č����Kr&�cً���>Ӻ�f+�}?k�|��� 6��\�����qw��Ĵ=�w���/s_2�s���5�$dVn��uB�|81 �"��$�/=Ol7����b�+�*�|ty�u�ZbϏ�C�]BN6���|�����c��Z����`���K��y��+i�?B��i=1�/����ܢ��0�ls�� ���N��Z�r4z% (����yb�;��;��H�XW�K�LۗՋ�QV�\�����[
]P2����`�E�[��6�T����]��-����<�%����fj�������}��/^n�p*s�S?���}s��X��O���g)�����*D�N��0��L5���=񃊟�����/�U��f�ﾋ��Ļ}��,ۍ_V�1E]�|��<�e����Mz���pS�P̯���+��۰̚	7��W��	�`Z�cco�39��֐u᝟��Ƨ��/�_���@j#o䖼#mn�]��k[��rEW�坱;A�6����"���={@Uǣ�m�,�I[r�C�Nou�(�NplA�ڿ��2�rԩ�=wF��?�t��N[x���I�%�|</���o��B[`������<}Dj��m��_�vTrd�:����BN��Jur_�g�
:�+!�#�6��@��;٣J;|�k�.�g�2�����(V�*䬮����K�B�ǩq�^x��:Vv��(]����R�g��ރ�R�_���jEp��{��u_��F�v,���zQh������,����v�t7��v�e�v�|���E*$�5���Jl%�ێ4Ҕ��j����i�l]%ĸ)�}�� Y���$�]�c��|��t~�`v�c�7�YAG�#b���hR��:D��2z�����:�J�]�߈���F��#j7�����R�I�7!�>z恴�y+��#	�["!�?�&�e����w�O~U2��&���*qq⌛r3כC��t���x�]Ϭ+j���C�S�H�G�� OdO-����kA�* ���dj�E�{}���c����g����h`*g�}�c���n�����3{F����n�f���C�&�z�+�:���WX����Өo�Y��Y���}��T|u�y �J�L9��#H�C�l���_>�./�1�&���O�o�����b�����ׄ��o����o���õW%R#��KOs���uOH%�x���.<��ѰB�v}�E����fT�i%O}���fL59gntr�rvԉ���q�tM��EB�8	T3��_�mN�A}Շ�4T��=�)GŽϥb�HN���@sQ�Yu7�k��g��õ�(%�7Ӱl��������$
�w�|�Q�[���)l�揖�,�󺰺�""�A��<�(-e<�W����1� ��1��V�`*�{N;�bC�e�(L��}�S�	�C ����f)�;1�1��zKX��>��B���-��"����X��W(w!z뗬��PÉa*Cq�'�U�̆ͷ?Z��m!W����0������D��3���<����a�,�p���d�}�4�Wv;F���k�#1�`����_4~��f.����9���:�d�E"���֡�t �<��mܟ��><4�m�����`L�Ώ�I �w����9�Э�i��^j���#��ì�����Ժ�G�WH���M֯�>[t���E%��3�Dk_�x��z^d_{��C�:$^�~�4��=�|Ԃq� ���~�"��P�%�1�ENȆ��c�᦬����k땪N��-}��i<$����69&��@�̨w�t�y����Vm1�n8��D��u�4�'Z�=��W�m�ާZ�Q��zТ�7����j@�T!�<ƾbU��b�_,��x�.6޶���/@>�>�	��5zn����ѐ�:I����W��)y�����:��nޏ.hl�RTZ��5x�V��擃���)�����G��>i����צ��گ_ W8�g��X|]�,=˓Q�rܖ��&���㏮y^���q�Q��=�{@�5�k������u@�����u=,Kç+��u	7�tF0{9&����@�YK5�~t�/���4��������z��ͺ���a?���n3>I��+Ժ�77A}��f�$z,Y���.�8�c�uEr��3�3�.��W���K�H�.���g]Ǹ� ���N�Zبa�/I7?�F9W�G��7>��FL}�yL�-4z8��	�����3z�b�b`�NVQ'�B�r��/� -��f[fCN� (�f�=]⡃�=@���r�.%�Pг�#��r�^�i�k0���O�;���Gs���0�ĝ�U-$(��޳�B&���@[��֎6�p/<d�߂tR=���+ߖt2#XXj~.L�$�`��w
��vamQ�o3�_��6�籈ͯt�T�/#�s�:[]Ķ���.�����W���?����4;�>��ML*<����^C�!0�d��'���?�(5C?�����5T��>�,5g���{�f|<JWBThc�*VM/��T��	�����Ғ�6��@�r���7hk�C�m-�d!�UҧwA8�ڑakZ�ʅ?�j��3�]��NT6�p�QW��	:O�_��_>��]a���J ��v�
 ������4s~Nϱo5�t��0���޿��g2��M���5X<�9�9g|~ɂu���3,E�~`)���Z��Cg8�|��d���3WC�YZ�s`��_db����"���ѓ���@��!�[�y��,�n���"���n��>h�;��r���C��;��{�ǲ>�W6o�\�w��~������Ն������@��ܺ���Tt��4���l�vzpLد���G$��v�o��O2u��-H�uO������iY����X��i|W��ڗ7����3���F��z�˜bbi?P�yŁ/m��)_����^l�䬽�a"B�/v�Kl1&���?�F�^��L�~OxXE�_k��:A�����Z�D��"�U#[<P,E��-K���Y�.74b����Y���]k�ET�/qa�
 B��6�K�4PgA��]�����me�^���J
��mA�:G)���.���K�։A�}!�9I. .���zY����ʬ��-��w�Y�=�t|O�/�즫�q���½��j���LǯsZ��,��9��&��릹��Fj�^m�^��P[��ĭ�[DKY]$��O�\F,����S\Bf��Z{����.NV��p��Ȣ�hE�-����>��������3�NORa�n*+�J���!��c/�a(1�᫑]ηc��f ��ԑ�}ƕ����|��R[v2�3�m���Z�Ȉ���+����z���y���v+���IWw�YgqS~�d�"��C�пƮ�qz���\������G����ܪQ�g<"�
���u�|�g��j}����x�P�{u�;W8����_c�ĥ�r)~���ѡ���F�(0���\z�n�ןwY�jC5�|i-(���%��;(*)�~�<�VzHrc�n���C��	��3:u�i�8������L�@�ی��ޗ��o��m� ƌ�=����%yh���-���z�7\��yJ���w�"¸��+N?�<9���0�Ѯ�>�]Vr2��C-XHVܾ�����_c�I��0O���7���ɴ�â�[�gV{{A�_�}��o���5+
�LuV�%.:I�D�+�Ykٗ���C�ִycE��������A��)'�|�u�Ӽ�n^�%/��@i�w��Q�Z�uO�P��]���n��A9O��ߟ�{��m�A��)�Nz����+�S�	��|�B�4�!]
��f9,��ѵ��\��#PR���[s������yz5@�@A�2�=��z�ǭ��m,x�ߎg�,̐}M��+���pk�\�z�Ao��.J��@����1O1��ۏ�4����.���Ɉ�ȵ�ư����J.i�Wq{�־��{�m%ag���S�LFQ]��u��B��b��6�X[��������8�U����:�I��fe��zv-��"͒u:4�p���'����&�Ѯ'66�j��=�űZ�Oj�����X�Nw���K%� %�!�ي��l���R۵������:8]?��oEK��I���Ҩ�ߵvL��#�W��AV�B�'0��ε�!�{� ��{�b�#z
�zZLk�
��*�M��KE�)�)�+�)�9�Y�+%�癸F�'����Qߺ1�7��L�,t �ǆC��Ww(;��勧v�K�;�Kj$���Q�p����	�����޵��A�~	]��3���h�V�B*�M5�,(mv���H��΍�~!m�4��h��0�v���UaPiCcOg�u&2�>��U�9�.ї�����_��Cǌ����/���<���+�"p�p�CHe#�a�E#��cd�S�!�w����d$�S=��qW&���Cbi�\/�c��K��Q�*�z����Rk1������*To���G�s�����u������������Z�Aa���^`�fS2]D�}w�V�4��efL5��K�6�4�M�ߊҊ^B�Z���}���M��>�=��Oj5���?��z�ձ���Hhr̓��(��b��m�uO���L�v�l�F9�D�P����/�N6 +8ѷ�(c�Ua�')����"��E�֤٪[����F2L�P3"�rz��Oަ�$��C�?��)Īm��Ӱ��	n�Ky�<]�to����ujƱ�S���_o*s���W�=	ߴ,��=|C����}N�� b�N|�!��C�*��)�5�ݓ�-��~̉D'/9;s�<��3��%�v��=>���x^�����0����>{�[���[�o�ؿ�0�<�LǤ�F]�1�SCF�<�z�NkrK�B�SYL�E�s.�3�u%.�Qi�5� -����Q�3�dK���{g=gRc9a�N�*�a�uM�J��o�^=ĝx>�|��}��'ҋ�#������R�����;<<C���/�*-B��i;e���u�޺�ٳ:��kZ5c�+��^*M������P5<�v��8��\Z��.���d�U^oU��[�k$"�f�)������wS(��*�4���(�Y��K3C��&�C�+�`���ץ쇯F&���Ґ�h3������	�ɝ[���I�D���F�����j�$@9��lm�-�|�c�SO'�����?Ӑ�^�aWUF�����!�d����.]�&QG�Į�Us�D�^f]���tG�s����g�p!��-�8}-�:޳�-�X[�g#�vp��yO��=�J1?ߴ�AE��:�D���;�Ң���LI��͑��{���t��2��@�7���ġ���e.E��G#`<�r���է�5�\/GKn��X6J"^&}��O�}��'?��<�Z��ɘ&��M�ӿZN������?��x�mgA���Pc-㤙�K龲�����W�`-@)u�R�G?��:e���s�6p|�J���<4Jʃ��f�v5��V
]�B��A}٨!�z���ؠ>i�t^ɟ =����<��`@��n{2��KŊ>������g�x�� �	�Gw�_^�l��]����G�GFp:�x����7J뭭4��(Ӳ����bf������(p��L5���b_�����rlio�S� ��i(�@�чu �޼���Y�/���k�3��N�v�gn.ZVp>]H G��Ɛ��g�p�c��$jY��mYf�l�@�����Z���L�c��p�%�d_ŋ��i�0b�H_}F�9��|�#�F�R�*5f��ÒnzXj��+�g�
�Q�p�g^FV��DK�8������/6^����<Y���I?JG�뛘�����f�nQk�P%�lY0IC�JJJ[��LuE�g�e\�e�"@w��w<;A�R~�)�a�����b�<�D]�����a��Е��:�4z3�Ώ�D}��V��~�p� �?8�2 ��ZM���[Қ\�0|a�jɵ��a�zI���C-3r���Ϯ�jk?��>[��(��ҷvo�hQ������OȬ*�ŢVf�<@֕�M*�����E�I<{\��f_��W\��R�#x_[`�
¶ڜ&�0]�ѵ=�ɯ'���p�@W�0��xR�v�v���pY���"�/�B�ѣG6�qΜ�~�T<td�R���+��;{?�:��~�fC��w4�"��� ��Ɓt6<ety`��QҊg��
�(g���]C��{T��\f4T[����-�PrUBG#B��_}���b�Z8�a�1�iu�Z�b��!C�TiUl�4���%ٕ��0��W˙�r���&��oc1n	��R?
�mP]`z]������E9��*L:��peM���Xӯ)Ġ�*�^0�̞>U.u�(ƕ��]��"UHeL[��Mx�-`����&��/ �?���L���H#ZC�}L��-a\u�cx[�Fr>����B,��NYIQ�k�����?�4������4���JKB3���p"�0��hই�a�.��t\�#Z;�g�V��m��-��>׈��OA�}��48�d��W�&��Xc'��6z���b<^�d�S�<Nf�c:^�8�$��O[��'<��%vxq�s�a{�� D�b��/���2ɣF5�a(7w�U�zJ�������9V]j�*�ui��d�#��=�@��<V2�p]ҫu���
��R�i�����-�"mX�)]�[���^D������
6�Ɲܘ����et��p_�e��'�^'ЍX��䛿���Kk�`"�G([�\�Ń���-%�b�a�Tsz|��}K>�*ܼ\�ه��3NZ���P��|c��L50����|��\�9Ù�I�(��̈�$��O�dВ�''�6$����Q�ۢ�:�a[�`������Y!oFT
;��,@_�U���r����	����<��2��$�5k�m(Yφ���E;�a��O�YҞ}��r����`	�]R��I��60H��}ڞ����E��\��+�B�z��4���?��{��=����?`��~�H�o��r��IT�2�"�x���o2��>gp\7���p'Lo�G������c�~!��no�BG@,x������9{����k�@���όB��^z�����,�t9�'`�ӏ7 e��躸_��=I,a��.q5
��m����W�>�b��q<4��[׮ǣ��?J$�T���=�vw߿��?�'U&�2�MN@��RzL*�L���u=fE��WM���,�O���5�4g6ǽ.u7YG�����G�Bm[1��Pmbᑚ������~��a�8>:�B���TV���Iy��X�Y����=B	J��1|DV����cv�X�ϸKW1%�T6���o�V�c�V
���şo����n��)$�0��L;�5Y�չm�����?H�0��<P���|� �@���`�,�Έ�kQpV����S�f��:�6�k��<�Mh�V&������~.}������g�ÂA8.�v����Ʉx2���^ڭ���8S�>1xA�����.䁷����#XPP�+g��L��:��o��������L����/��~M��J��$�����_F�E�30G��8\�H��6�����Y�L��o�il|D��D��5���F��bf�F���G��9D��D��EE��0q�W��F��V>B;q�Lꭔ��_��澋��>�ܮ>���q�A��C*O^1��ƌ=���BG{O�N�|;B�t�m�?�����Hd��;�.f�"F/�����6��36��P]�&���4UK �<��$��89v�����jWv��AP��!1ß��Ҿ�F�}�ٹ��%&�a�g1����vl����#��<�i��]{�5wP���i���ΌMy�:W��k?R]0��A ���W!�6���G.�������Z����S�~�ao��pm�
{Ķ��I9{:�������0���C�>~�}�F�Hj�G����aj�� n��ԩ�C�=��l���Xr����ݙC���_�$^�t�5�G|�.��&�~�UJ �hXym�WU����6�ھ�Q��t���!�v` K#]�9Y��?�YK�Ÿ��3��Q2¼5��s�#fuj�-��U�x�}wd��5S���L�����}`+k�#q9��%�4l"�A+�_`���gLq��z]�����I�����g5'&@�|gwm�2"�>O���bpN]����N�72Q�'�)\p�io�L�}�//{cl��gc����|�p��[�)��˰㢅ؕ'Ӈ��X�FCiM�^��qm�'��U۬��'��4��Y�̜�+R��n	��
d�V�g�Wd+kE,�X�(�4�/�,ؾ��E�S+�n�6����8FJ%𚄕nw���g�UG�+m��Y�-R�]�>�x�oOȆvUa��ۘ׵`mh�.@]���2���7�]��O��`�"���֕6SU#�#��KG��o+}@��z=���	�u�K���∯m�V
A���B CQj^؋>Q�;�cnޅ����|�����C3�Pa�~pf�ϸ�=iZ�I��\����ܱ�Bk�ugq��I�J���?�z���U]�������毕�!=[٩!�֝��S7y)�� Ĭ'M�����$1��@N�}����|ˍ {7��ނ�>��%{/���$r��Ͱ��5��tD(L��?:=#�����ZF�яred�o����N�,fk�o�E��bq��9Qσԋyh�z5�w�n"����P�k)���2\Q�..�a$u���:��-��S�Q!�J�����%޽���|?��,W߼���S��+���;��1iR6���Q����G몆�C��#���\��G�Dh!W�`���j��o\&�o8�J\Q�H���ѦuYI'30��C�j�1w+���ܒ_��Ln����f�jg�<g�l�
����~�]4���7�e��7ڲ=���\�FE����`�OՂ��m<_��;����u���^�H=��z��q醧�W߹��k��L�����Z�\�ۮBC���46?�EС���A�K<"nk'��T�M�dz�	�r��,tf��ʫYf
jR~|O�O>�m�e:���g�,X�� �g����	�M���ݖ#���������2�^*�h-.�����[d��^[�;jX6�$�;�Ղ[�b���˓1�u���������[� �h�z`�*s�w�)\�����T�p�@H(�S���:X"�k��o�Ao����H[�\��lC�5����<�D�q0���`�/'ei墺�������c`5<�;q+|ǤX��I��3%� ����Xu+��J�>ås��ow�M����~���D�V����i"�]���YDw4BE�6���z���Ju��J��N��t�(�b��C�W;�R�
���"J��������3c����F(���@���YAٻ�EP��C9�8~�ݠ�	��� ��ڜ�Û��ӈ��������9"Y$=�����:ɢ�Z��}��+A8��m)�T*�����>f��1�g��?��/F��=;[�K��:ԓW���Ⱦ�BY�T!�a}@��ز��ܙ��Q�<UćXix"���SPZ�}�^ϵm�/���3�p���4�T�[;�S��̸�b���>�޽=�;��W!d$Kᘤ�)o�����f���1=
C׫��Y����U˯MY�Sf`���y{gỚ����r���4���oߓvKz���<��q����r�KI/�^��U�!����ᘍ�N�������$R��`U�"V��f��;��%��%&��^8k_�T�^뽠,��* l� _�-��(S6��`x����H�ߢ?_�s������Kܝ��ޘQ'���ߙ��j�����:�e�20.�z�.��j=�%����YE�G�O�s��g����>JV��4�F�z���"C��X�())���2�2?�愻�GO)���&)=ֶd�@҃��qy��Y�!C�Zz�T	�zt��v��ux�r= ��`���|�)�ߘ�Ŵ������ʩ�{`��n;i�f�H��;{�E�3��s{Z�f��'Ԁ��y�H�,����z�/��T�VU�R�iCm2|a|�<��s��̓{>�u��|H4�=�G��-4�Q��'�t��ըO	�'N�
����~:�`F�8^cB�>�2E`�o%|�hkjj��ּ����M�*����6hBWlw�90��x4<6��r)�f2$�:\Ig�"*�V�����^��L�1|�K���}�͆ڤV5q����.K'S^!���f{�*�Yh���*:+j�3g�Xhrg�&�,��/� �L�פ0�-�!B�>�JR�	�6�HWh���\ah]�*0:������),����-���Z
������8֟c�N�<��w�k�Y�\�G�~��k�:�|�@���|^kcr�i���e�Gz����Pڏl7�f� ��fu�>V�si=��z�<�����i���?қH�E �d�����c���;��Au���+s��*���>������m�������ΰ4������#�l�|&��ǫ��zA}6U!��9g\�s����W����Iom&|���@$��`���V�୔O�ki����0)��w���1��g����ݳQ��`���&B��1Wֶ)1a�:;?,���Y���V�Y
$��.y:%����#�,���pɆ�@�b
wd@H���Y��؝���L�eͳ�O���]�^�*��Z1�^b�$Ϝ����Y�Ay 2�y*d�C�����T�(05�[��C'��Ů� 
�+�I��w���%�Ũ�=>���&TH�
���Ћ�����;	�{Ք�'��k�1�i����r�N����XJiD�����p��W�����_��Hb�3?��?7�m��e��T�f���Ү��݇B�/�g�pR&k9���6z��Y:��q�[��~��)��|ݠCD�g�T�P�}*�x6������_uf#yR��7���u��x��M�%�'�Ւ��b��:DQ���Ve�B��O�N+�4�jx�:/�Q����;��J���<����ԃ5^cߥ��=�W|���2�����u%�����u���7
Ʃ���V<�>\!AɅ)�3:��q��'�C�A��#��e_Ę�{���Ʊ��� ͖i��5�D�Am�k� ,�Fw����
WVl)��|; 1��>a1���
Y�++�]�@�{�T�~�����3=��لz��V甽-	������n=�����s�e��f�*�=*��Ȫ�S�jѯ����c�P����>�=�E���sy��=�7���CL�8��C��ә,��0�fWr�ԌI����_O���R�qp/��逖N����������A�)i����ӥ����/DP�����,��J�����R7	 �6���V�!�5'G��3A���tgW����a.y�Td�ݱ�Z**�vA� �W�Q��jR:��֮Y��o#x�6,�A��x �۵����XJ{;%��B+oi�~	s��Q�qj2��?d�xk�~���`���I�P:N.�������샸a\�Tm"ݟс���W��/�j�b|&��3����+�ߞ;R[�J�����"�\z���'�����p����΂�$	L+*X�+LR��M�D�y���}r����oe�;�z?��"���iH�Tu��D���r��dd��$��%���%㷶�'xy~$���[L��/��`�_F�������o�-9���2>\UCm��S��P$���Ϳ�0Aljkk�%�[f�n�kM�`�@�w�DO�� G��Re!b]�}�{�n��#�n(%x��� �do�vj�
۬cC�V8s9�5����hU���':J�z;?�/ o�^I�,\x��6^��cĮؔ��_Ot����|S������RT�Aꉊ6H��V��
�KO�Ԙ f�o+�c��z=`�~8���?��䩮��گ���è���Rw�c͔U�أ�2F��#��o\�(}m�7����>�������,�;���ط�䖤/��,��v\Ȩ����䰿�5��kba�@&���^f���ӮDŏ�y��Q)m�<��ۧ�O��0Y�40�<�ths=����c�\K|vzv��oK>��h	5T������޼J�8^�R�(aff��~T��1e�Z�D��A�s�Cot��"iSC�����>����8����W���*�7T�  �-�^������M�4����t�y����ܚ<B#ڄ�dd���xi�R�z� ��y�P�4ܟ;�I74���Ȯ�]~K�U�=�h>8�怡�v��/���əxO2*Mw0���.�X�5���7fx�g��<����.�q	��O���8��*A�Wl����_U�h�i(��B���шE�2t��jz2S��N�s
�z�{��ɠh�;t~�˹�ó#�&v��>{K!�ye�O��"���ς3�΃���C8%:5�(�������1���ʠ�E��J�M <
�K�d(!����݉�ۿ��"�s��yFF�����	���M��k��ĺ_Gp���+��4N���k�AQ_QR��ߜ$3�K(��#@��X�g�5��[W졒̦�/W�9�����)u*yY'�>�����*84j��;Hz���z�0H&7#�;�9��#����Ku�\"�,�����kf2{�v/���uw��1-�4����Z[��Q�5t�P%)M{U9򦯼��:^̏�7Fq!M�\���#��m�E�I4��><��Q�1DT׿�Z��+LB���]����ߟ3���ir�ϔ�f����VO�on���9��}�D�79�/cz�p��8~��l��M��E� 5�|�%}y�'�-afԱ�!�K���~�cN+ZL�G���y�pV�=�(�,���N?R5����	?��,d��|�_��k�`����q++���j��O�ݯ�v�u�����cYp��B&�-�y�&�O�j:�=��'�os{+����3$t� ��-�Q�N� U�����K���M(~RV�L���
 $�*�����q�G9_;��A
�O)�uڀ+�M,�·l��>Z�ض�RY�Vw4y�7� 1��Y���>���M@�8LY�u�y���А��RR.��k���| �ٮ�(������e�D�nO�H��_k��=t�]�^����銎즾'�o%'��c��Yy�f����fZ�bD��.)5���я���"�����c�!�=`�m?������H�|�ݵI���<��4#���������(?����F���~���Pq��<ᇇԮ�x\x�|z�'��w���f��X^��|�+�P�{�Lt?|���j�T�(҉�|�|�|��o�|�9�َ������t7���{�W��`�]���L�P~��9�!�+P:<�����Zc ��v�Ҫ�nzEP��oۿYa��3��_�=iC7�>_2��@xlHד������DP�v�w�B:��wj�w����9W�����L� ���e�>����_b���{a��1a�o��$ϟE\���j��_����s�*������,[�����[�`s/�d��z�Uִ��5����|>�3���z�v���j�����*��*mӆ�P^���9���?��~[�k�,�Tĕ����x��$��?�
\y�yz��
)��I'y�Zg [��Lu;����gv�������u�:�2��:��(��lݩ%{��������"y��y�C��uȶ���H�
����֌9�-�JDr���:���M~�f�|��
�y
�1|�oqE4zC!^܊C9��d���2����t�'��,c����`���ȁ�q�'[�I+]���[ь��<`!/��f�0//_Y[�����?�����͂�{����;��|#(  ����TCY	'�bؤ�ζT�_O`�^�_ZC���v�e�(�e6���.��5��Ў��a�;}��<;|�7�ഹ@=���[{k�ߗ��-BZ<VV��������Iy�\כ�<��t�ft.�����(W���Q�W���%��akS�`���9�����@�Ǧ��OA��lk"?m�zR��Ow�d_�J��X�I��s�>����_�nw���(u�	����"n�?��3���Q{� ����ZAZ4vjTl����{ﭤf�E�Y[�;�VI��YZT����\���w���s߯r}�$Ī�s�fu�M9����1E��q�L��F1T��~7:��� ��2az��>�/��/3B��zm�dPZ�\Xh=��X�q�`���*��8XmK��s�������NDW�u �=S�Ჭy�}FE8 �A�_|���i�F����׶d�[%I��r׍��+�cD���uO�t���-HJ���d2*)�j_��xf��:�F��f"*NĿAW?K�w�o�R�ߣG�;)�vѰލJ
�p��>��|�-�x�y�.Wǟ��n��8��,��\7��ū��u���b�R5��I:KsC�]"�I:皝�W\ӟ��:�j�q��X��1<b,�_��ܛ�z���'�����y&E	�Mw�6��)�Ylzx������
�'vQK�ٯ �'���)�"���t!��U+.�.�s�U�C���*<�6ö�Z����<XO�I�ϯ��3���^-З$H��1�Y
�E`�0� b��I^�d���R�N�A��722s�z�\AY��ǃ�0 �t�Wd�*��3�㺳�5��Xn�Ej�e$
P�)!�dؓ=�~��򜷣!�:�n(6�����^��YC���!��ό����4-����e�_���'��8�;z���{����� ��8������H��2���x����H�����2->���X30�cPf'�d�cj�V��$�Y&��ch ��#v�����=0uy��>�1"�̧�?d@�}�B���B��o�L��I�UKw/��ap�"�W�V�X	���/ � ڏ�a�J,twa�L�1X}V{n���� �4�W6=փ஍^��Mɠm_#�zV�I%6��ٲu�Zr��SM��3X5�ށ��������e����.1h�i�V}Cfv����g�<�%m���C~���w+��3j�h�m,9oK��fY��E5��ՠ�m*|�����愣�r�sdV���@J
�W�g���b���T~4���0����9��Ud�O��P�& �|�`� �(b��*�3ɂx]��oS`ʊ*kAS�~����k����D��� @g��&���
=�}�&=�}J��Wm��G�b~�ǵ���;���0ޓO ���w�=������c�+�|f��~K*H�ܕ���4��l�;q6Ա��~��*����I߿08�vѰ�#��}����9W*�A�B��3
yn��Rx����Ձ)l�����������Fi�*�$ ��r�%Q�������F��]%�|_�jVk�.�_| �P��/�>ܯ���n�F��y�$=mT|�����������?��� �l��~{\rhN6=�D.6�%�����~E�S�H���|l���{�#|�����w$F;r~��x#�y�B�F*Z�,�o(Bx���9�ٵ��m�����)�l)��%�cV:�՟�����6!�8���pU&����>>�"���:�~�>��IS՜ �`���Z��J{��p������ޭ��Fj�9J�"a�P��<�/Z����@��A�������X�eoz����xi�6S1ql�~�8W����N0�+X6�A�/KzXBvf1=��ä�
��`��/K�bq��r,�R�1�U���G���lSZ+Zcծt'�wͪ`$G�����Hʇ7	�i��MM��86v��^C�[�~"��0lz�	�0;
����X8��o��ආ�4TE�#N����ȳ G+ɪ6���A��L�
?��?uTc-��1O<Ơ��ci�Y��9�ԉ��H�29���Cq���Xz�q6�ǲ`����c��>+�R�љ�i���Ɯ��Ձ��P�ԥ�݃Ο����S�dM�&|��	I�`ٯ�cʰy/�oX*�ͺd���F,�HI��ڳ9�Ѕ$�X`P��)�*|;� �_!sڈY�C�����Vc[��C��54����A�i. 7:�%����.��-j䍨����E���d ��6�^1�Rf7W�4������ЊCm� �j�P�O���{�Xb��HHeɧ����RZ�؀�US�J��`y| CC;�Dc��S@��s��C�L�P�Xl�;i���	�)޻���.Z(�E���/5��b���"I" �P��W�qa<2Ԁ��w��h���0�U`;��+,)��xe���R��-�:�ɩ���)���!���[eddԝ8nĬ�k0�%2>ֶ�º��}e���g0�xKuk�q�ܓY�d��*�
��f�ï�������KսH��@�"�ǽqF�g���;���_�\����]~���|1ɟc��0�������d���&�_�R��=��a�dKz�p�nvU?�bL���์/�0��;F�_��B黃Ot��3���,<��9�W�ؤ�bB&���m?�����[�)N�2�.��[gC���}�Y��[�!"Eܷ�e ��H�j:pKG�z/QAu�'w^�)������;��ۤ�S����н�~�����s��3�%�L�Y�!VY��\8}�0�&7����L8JU������
��x�X�ٵHh��.m��I����y�Z�Cv�F�U�E.%���`)�,�Ƈ\4̿��;�_H҂�/2ۀBK0A��l���U��#X���~����01T����%��{�wT�D�\0�V�7��0ԣ{SR@����lԌ�}J���QK��>�ۄ7��f; N�C
��-m$�\%(+ 3{���s��.�*���D�X7W��B:M��i���C�'G���)t,�U�����xЉ<�Y�By���RŒ9c�Dǝ��������	���@5v�_lX�C�y�r.(�(mN#���=��q|�Yl0�#3��b�~�"�l~�}W������f��e����{(J�oka�}Cpjn�gߣ��D�ϐ�����|�z+V���cn�d��D�B�Z�gh2�&�^���'l��DPR]�s�q�S����T�ҌM��������{ ��7<kw7��H�p�ft��|����i�qP	��jό(^#S4v�bر�z��z6���%8>>�SbX�)�l^	Z��F��!��R5���gy���r=�R,?*b�<~����s O�����j�����ULF<r#>�,;�n]�n��{�?.�@"Sfw��\h++C5B�B
}�.����WI?i��^�ʠ���2�hƺ�I
���*e�o�փZ�|��Q�:=�Ѹ��=��V:;ylN�R<���oU�OH���C�
	��Da9�圎�ٰR����9����|�j�4�U�ޔ
f����i�����8�Z![��!EB�i�-x)�cċ��+�yk�� �Tm�x�4�'���*_���C �Lը���'{��g�}~ģ]2�aIl�t؝�41Hw�4����� ��������l�⊇l������?����ٯ����|x�������{�l��*��^�Dz����9��]��(��q��ڙ�Y�S^���3o���o���.���);]q/T4����\_�w��B�<�C?�~0_����E�������M�Z����ޢ�Q��>��1���d����C@�Y.�2�5�Np?@Q_�jG&�g��Ӗ�����l+Ơ�m�ȼ���Z�%CV��f�YI;�v�=Y��z0����װ��d����7a�ݔJ�B��l��Z2��P���}ԙ�+��T��o2*�/�R@pכ��k��}��5����Qe\����|��R(y��g2j����K+3��R-
�!	Fr�p�&���=ˏv�̰k�)��	���.)�)��h�Y��G� Ɨ\�o��1��>m�e��1�]3�+��[֮�W�툌�io���ߩ(�K_�����Rz/�]�0z�j�C����ʄX��T�n!zۼ1"6��7�;��~cv	W=A�/s�#+�M�{���7M�g����l�a�;�9��O��Z����y:Fq!D�>g`�3��C���CQ�<��o���p/�p�8��G����ퟵ�^4��-:z��"_�2f������@����DK����5�&qXAT�5�ڞw�"b�ǲ��E&�wM�P�9b����� ��6&I�I���0�y�V���7B�V��s���{�J�����P:+M͉ .�<풠�Y��:Y(g?��/LNZ|y���� �u>Y�o���ܽ�����a�0ô���8�6ΊI����CX��)7�O�$Vz�e���d�4�[�lJ$�u���V��3��k���)��K�&��s�>��d�O��ka�f� T�&��d��('������(N5�<+��{zӆ�P&+���1O
����L�!�c<��q��;�7�Z�&��5��7��1Vq�\cu�|(�'�aߙ7�t7���L �X;J*�G�JY��������Fb��8U3"gg���7V�Py �PH��`N8;rp�0>r���0X���vE��O���/r'���b�+��@-.�����=�eW�o�2Me�e�u񅾅�fF=��K2�ߏ[C�EqC%��M�+��p�7��>�1(�$��dH���gw�څu�_�Ђq��,Y�d쇯6�Պ42������Z��J�t;B�=��|�^ �{C>���_@�6�ϴ����V7��m	�̨�y!:�=�f� p�8yN���q�{K����g�.oX�T�����-a��V�eK�h�!n����S��Q4�x��AR�����3�PU�q�O�'-�(5�[	�׫�|��M�z����n?>��N��3��F(܎���aJD�¿��_wH��{�S���ݯS8����׌F�[d�1I��4�ӗ�|I��nc�8�u�2x�I�6�[VhP�����%����'5�Q_�����ھ�{Cfb��9{���V8z���8��k�<�!fE��)V�Di�7ڏ(ߕ���XAo:{����,�9`���
].��)�\��$?n�'��
 �g��R���o�S�]�ɡa�ه�2	���5��?#9iǬ���<}�wb&Ξ���[U�ť'?�edx��U����;��|���&*�����)����Q^�h��M[��&
9�ƛE��D�̭�w?����9�b�������Z�k���&6�'[�R.</Bv}�>�A j"�J�).<`����p}_D��+�|�f͉tPsi�^��_��4�Yك�K�D(��@i=�,�6!�D�� ���e�?[�ͼI�ҕۋ�����A0��Դ��n���S\�v���"��ż��x��i[>^|)�ہ緎�(��@��f���,Ϳ~�rc�Z;S_�=�z��( �-�\�7��~g�������<+0)��g�e<>���[|iQ���ʒZ��?�'���۪��M�u{��U�r~�Y��\QPa4�{�f�'s�&6>�h�פu�s?��	Aax�CϛzH�Cڰ��k�t��C=�b⮡��\��O�	VKG��1[=P=����R�71�u�.�yx����3/(D!�8\���M4Y�!��OT���˲=�>��Q{���xH���uЂ�CK����N�4��B��e���R�?{1���YsQ/�욄��*aЁm���x����T�!�w���_�z6kPKsN��J���sZ�7:*�bg?�5ȟD+	���N�E�n${-8糆K���Y��"4#�Ɲ�'��6�׎po5�$HC��L�,gY���{~�|A(cd�[ο�LXK��Ν�������i��X��J�ĄFF[�؎���%�JJ#�ٿ�

2Ɵ�Ve�P���	M.K53U�0J��l�t����4Åms�i��[����k<�n~t`w2m��������������ǜl[n�����-��N�Yl�P�ϸ���	�*�n�V�m�[�����H{r~�մm���C׿@5gE��{NֳG�Bo(Eǚ��ywk��c��θI�e�b@���\�N���%�&A��7*���Q�����;��V�6��	�;c���ܞMY���W�n�zæ!���O
E+)5�����+9_w��?:�o��>��݋Z�����P&�A�Э�M����É�k@��w��(�xx�ZM�U�w75��n��q�я>Vu�/�O����.
C�sk��-�9�&�<8)����) �'�֩貥	g���,���ޟ��$��nM�� �s�NlgjM.4�|�|����ȓ��|�uR 4\`G�s��gW�m?d<
��tu���^p^
>�Y�^<Q��B����D2q�a~
%6��M�O�Q|��|��o�FR�'2�<�@_=emЕ�O��
���e�k}����Z�����Q��e��P�5���෹��~��]�D�|?�������ϱ�9���k�0�Wn����
���Qt�}l!&}^s�S�dY�������.�������[�1�J˒��T���܍4'�gy;A�m�X=$�W8�'��R��5�ՃN{7o��!1����K!�e��'O�/sf���Y���tu��bkn�#YfE�D����e��Ii��f�C���W�>�����ur�wu|d����*��-��������_���3�smM�F7}=���'§��H`J�o`�LΘ��ߒD��������/��������5f"��x��MijL�}�|C����z�@|@�+�
S�P��"Aə�������x�
�ߠ�'4N;D�)��ާ�U�G3�-��\�����k�w���V�0���0,��S����M7�&��\�Ȏ��t8 	�����T�+��ЎЄ��&�ҭ�f��c)jsER��ő]2JݛƓ,��.B�v�XT,CA��aN���7n9�˿��Kg����h�v�u��9�Rj�@��6�H���aoM>yWb��R�@��.>����t�e�K��]�%_�W���5L�`V��J�x��w�/���rY�C�����|��'&Vw�\�NUC�B�χ&'K���pS�g�oe!�EDƱ\��S9>��@�7��B�����[�~~P�{�/O��;K�oV���p�G<�Z��
!w����N���s��軛n�+�
��!3��z M�ڷ9�lt%�Lyc'�ׂ��VˢsS]���K �y=��sˑ���"��:���E7��gi1	�8½*�V(�(�6�z�����?��_��!n��{K����6�-gЇϠ��`��2�s��>��\��Zq�|��cȓhL2�-��$�8�rw&S�z?��� 's*�N�q{�I���Zш��2���o����8��R}]6tͮ�`3oiz��qЧ$2���ɔ�7ͼ�P�)S���B�zH��#�NA��t+��4��D�n*SRY�	<��8d_�7�}>*���
�J��=r��'#��)�̽;oٺp��r�s�V�~��m�����;4v�;��McX���|�HI=�}� =_e�Z�YF�]F�����W3��u���2A�U�*�X+)�����A�g�6�nn��4�L����������Ҫ�Y� x/�З���c��z���,cL,[�_|����9*��Ӊ���P�n�1~���*q�蕙:����X3h���'�*{�J�.�Sr�l&�������{�	����bWi���~M���Pd�#˹{G���tF8̡���J�X�
�&�����t�K���Y2@�5髠Y|�D?���#�Ȼ�c�0g��E�h���01X�	B��a�q��E	1"��4�P�4uXE��Fj)Gk"̵*ry�zok��G.yB����Ļpr���=��X!���?X���A�//�BV��^�Y�RP����?�W��u'�Of�����gNZ���Lw	Ưط�W�/86w��^��l?�K����;�/)��S�'���}Wۏo��fǏԁW�Ok���y/���i�n����3P������){���P�H��,iBL�T}"4�z?� aa�N������l�p��WU�K4�-�L�/��a�U�=qDn����΀��eJ�5:�+�e��,�D�������!�Z"�'�A��.ۋ<��:������k��	0AH�t�U��,�s6�m0a,2�
(�X2��́K_�y$@�5>�ӶTM�H�͵�pp����ll�BF�q*���V���Y�����K0p%�(`��k*�(BM!����V��,��&"y�md�&���3�������;s�CB	����T��Ǎ*���/y1B�XNfA��rNR�es�dc9���̑%,�;f��!��I75c����;������ |����k�������Tr�����EaT�R����Ť���řQ�f�H��{�fݺ �h�:���R��_��/�;�W�K'�%�y�9�ƾO;w�����"��פA����M:H���l�	����=�U@��c��6�-ZWEv�S8]Z{"�2�E���Oe�CE	�]�_��]:����8�QA��=@�W� Z���g�ҵ�p���z���R��:��
�t�+��Hs�!1p8Y�s��r!��"L�_�y`�p�t�ؗ���1������$�8,����'5�����7D[0�˂� W³-G�T�PܛО��!��iކTEQ*W�m�l��TNñ�|~�CU�@F^�9�������9Ε�g>��f��Y�[Lik�f���c�k��4�Tk�c�{�:��'�0���u��&��;`�e���p
4MR8���t®VH
�#��(R,w��X���Ӯ��DZv��>*�d=C��/qrӳٔê��V̇/?嶲����庯-���ƹ[�����|���'�����41H����+���.��� �G{�R�R�����hW���ػ���h;9�A\5"�b�0A�t�����o>^zon��g9�>�o���5�|d+������9�%���8b������S����-o~Wix�֪Y,L+�`W��Oӎs��B��Ę�D޾jj ���Q\k��.�?f���zOS�P���p���W��)b�J�|���=����ZU�y�B'%��R�Kb�b�M|��uu�=3�0�t*��5@k�j^ �H��j(���4Dh��{u�$�sut�}���f7�����b��IRàC�t�2��]�����<W��3��a���Q��?C�ϵ&/V_��+���Qw�9����y4{uzU,�ᢧ9��H-!��P� �¿W�Z-U�q��koui�
����玬�y�!��B��1W�F!GWg�@Ucp3�����B�Ւ�����(C�%�_�G�W$���b�A��n�V90�4 �]Unz�&�5.|���Eѡx�js�v1;�8=5��Lhͬ�Q�/�&��	��尺{m0�6E�H�	]7x�vNq��d�n(���������t%�|ZA��r��.��)�eE��5����G�>T}�Mp�׉�rs^H�8�?��}��{]����SGZ&/��n����e��"9��.�s_�/�@�f}�i�b
�����l��U4��
��dh�%�"9/�l6Ã]Z��1���t��s�)�hz�2����:\�
��6Q�(elVT^3O�gf�$�r��-�����c�B��'Üb�xq�G

W�CV]<����T�O���j�'�2Oٛ0jw�zp���t��}��䄋���{��r}�Si�򜅮m�����R�*g�8�щ�gA�pޫ��q��W�q�8��;{��&M��w����{�P�����ז�4�r�~��I�W��)HB�j�6Z,ġ�<�|��q�������x��V5�5iKy�.��b=�a	N����O@���~�?v6Y l�'���*�Ao[L|L�keK�ւ�mְ�s䊾����H9Q���Mk�'6��h���] 8_�A�eP�yD��ľ�����¦Kj�}x�����UwSɤ���s{�,�a]�!qF�����nn����t0�|�Z�gHx���(R�w�'H�>!o|ȺG�@)p[/���]^.au�rߡ�wb�����������ĥ���������KG��l���^o�X�Y��=&��!������泷�����{F?ˎ[.r20�F<\���w�n?����:���߳!�4�� ����#�~��;~�Ѽn�x�kW���I�@p�x���r��[e7�����e>��崊�����q"h�YڄϬ��dȞ�׺06���q[:6ܻQS���37���}d�BO��d
�����Kӈ���c��d��^T��4aiӇ����Չ��� �9��*0 �����d�����hͣ,�z���y�z�/����*��\}z�87�J�X@�p�8��ю2c�)X3�~��� �B,2)M<>�p4�r�����y���٘�]N�]Y?�Lle9��m�0Kҫ�T�;nk>�c�*#�����.�hv��R����&�a�d�e����	��Cޛ����忞��E�b�Q��2:��:rj�	�Lh�z���p�[�0��;A�m�4��U@�_}>�U�1���;BZ��[m����Y�{�3~���u�z�e��O��g�׌�����{2BI�MX��w�⃹#�A��!Wĥ˿����<eF�0����ۅ@]d7jQ(�����j�|I�r_WM>9�υK
"���y�_+'�q�%2�����#���Ƶ���������`i��!i"�S0�z�;����{��p��I�
 u�����v���H�t��n�d�]��	 Gς�^߮{��p#s���k����ʸ2���"��UD7γ��V1^j��>vlo�i��&��h=�F��ZH��2�F�Q�����/�ήY
��� �KHZ��j�;�p�&6��
ԝ���W�}rkӬ�~k�,
	O��S�S�)]7����w@�C�8�����ظǟ:T�P1w����X��݅�e���5��2^��y����D�+)�L'?���KG?
���l\;�����-lDz����"��W��Z�����n4�;$��Pthz�I���������ː���o���xq�+d���mm�r�iecQ���2��6�K8*!S�WQZ�1X��
��E�[����ľ2����f�i��S��/yC#��2[����n�h�o0�e�9���ìz&$�DG�4I��nw0%Vm���ås�C�d�����5����$ԍ��� �g�`Q7�i~�3'_^A��s[�v��P���F�kP]5C�����U,ȯe����c����l��0W��w����(�N����q\<��f%���yOZ[;��嚂( F��vR9c�Z�0l$G@9т�-��-���
᯻�%k��Cm�u��_TD����o'��i���Qh$�����{ennNn�|�(W�N���:7=�F�o��5{u�¾22X��S�I��-�HF{�u5�V��^��'a�g��fdyca� ,����Q�`�&'������C$��g���#�B_J(�s�=x=���r�|:���)����d�T������-~�%#x�ZJ���П=��2C�����Zջ3�lޥ����:S���%]~HnŤdޛ�T+X�O�}�^�$��q�]2`�hɳA�ԡ\�׶/X"��D �3^�mnm�
�,Ȫ2
b�K��K�U�C)UH,a���BQ&�������p,�X��/�Y9d\�*��s}�z_5���魡	����؍�I9^��?0� M����*&����|���%�U�X������5�v�!D�"a	�L� 3p�>`�Ӫ;�#�!�hF�5��[w𴲂�����~2q�<%_����U��1(�*�����8�qy��N�[c��H���c�N3g)i�(��[S�ڂ�IV+�C�X����+m���0�|��:����L�T߬�1��U���ao���B#I�e�ϯ`ō����3E��t�?˪ah���w5��Ci�U�W����ۿ����9���z
Q0�[�������n2�.		QKq��Ӝ�?.������4�O%��2��K�T빋�mVX�i+hɣ���L����Ȕ�y��@�m��f�������>1�%�������UGG]����4�E(6��՛ۏդ�JSyz��
�+ݗ�3���,�[.W[:g��*wΑ��ty����y���1���NC)�>0�p%2f��"���y���� oZ�yy;[Z25ma���p��l�ʏOj�}�8 ~z.�<<�Q�[�Pk���#Sh�L�QW��O��Zy����5��h�������~��΋�˱��:����2-�����G����6R�.��8"C��>�W�wzb�g4o]���lZZTh�b��C�<�Q(���a�G��ꙛ�������v��
�5�����'Y�u��#�1�E8�C�^@YykYYd��^>�cs.%���݈�{����Qo�ZN�C� ���ڋ��^��^�a�,%�ak�T��H��{ވ��΀����1���H1A;�A�d�L��v�@��Nc����6N��m���س��M�;&U��B��Ⓑ�+1+�ex�V�޽_4#��h�W{��t6���Uڒ���u�Y55�^��m/b=R�g3��c>�]�ߑ�ї�7�o�˱ ��w�<�v�%ͼ0��T��m�v`V���������'D��f�ZjX�s�_h@�5+*ğ�z۔�HN�P�?�|;��������x;��)��R���j��k=�`�.ӆr;��j��`jE�k���K�%t�/�[H�c!Q|\��;�� 5��b���~��^ /��	��w̦5K��E5�#5.9=�B��b^��ҵG�]pX��Kϕ���l��������z��Jz�7?�<�j+��j�k*��h?��<	�HFH}�hv��m�e~q���u95�8_�B���Ht��z�N��9����XM$d������d������_��4���a&VR7�p����l������t���@΋�l��0ӽ��Yy���Z��j��0�Y[��"_Pu�ᐱ�=�p�20hXt������Ah�
�;��җ������&�ߑ=���iMJ���m��%�C(�2-�-�6}�>�u*�K�� W7���6�	���x��i7�ѭ�z{�9�v8Ϳ'4��mV��!�]���Y����B=C�d������!8	��Ⱦ�u�!�jg���P���1��9��%E���VDD�f3��Ƌ�61��߾�����^ŋ�,�V�%침5u�'�����E��ҳ�.�[C��N��D4�� ���Zk���ϟHGbr�?弽f�z��TDqbD�ƈ����K=�-H�8���vL�޸��D"u���1�oTo����-
֑�޻$pz�QtME�V5�F��9m�>wy�����\~�g�*Q�ah;Q�/����?a��6�����6����F�����out2�S E�7,�/�'�<�ੌ_�SYm�dZj��Z����!�쟁G��N�3�U�++S���A �ؿ7���h�f�ۖ�4�������'�`�\����t�S�
2
��v���sRۗ���{���5	�Eh��ch��ԯ�w̰�P�?�U�����`Y�e�I��K�^�N���cL0emM�}�{��AZQ��1��d���^8ґ�s:���ߦ��6����������#�G���~-}af&F`N�_�~� �%I�̃�`��o�a�!�go�&%�@�fd�5?�����/�Ȕ)hTZ,�R<K?�����+Z�Գ���N�U�xk57^� iUfHGKh����+�6�-2-�Z�w���(*���|������C��+�h4���[�
z�jHWm�kC��!Y�
��뻘8>���a�}�;�@�0�9��^��w�go^�I�ng�8��ɣ�_�S���}(ޜ�hs�u`?�@���b�hnw��`�d��|v�ֆ&����]���R��Z}���~G{��C3���">8��
�c��4������;1�K0o�K��r��]�1���Ϧ�,~3A<��^���^��fGlb/	��u�q@�۔i~���*�4}|�r�Lǽ���ߣi�E߃��M.^N���g����w���t2 fؼ�b֞AS��'��W}�W�G>���;~`��uh&��	t����F>�2FZ�?U��-<�8M/|�0�Q���'e*��;����j<�h�]���RLy�NLL���ބ��꽜m��zp�\�X ;���+���AE��J5ԉ&]�Mw��qJlbz�{��~����(�����Ń ��B� >��
M���C�_�x�v���fı<�ZoOi�Q����+և�N#�
�������������8��<��Ih�%���OP���n�{�y��@,�Z:�!���yB��7�4]2��V�p0Ԇ�=��6U�	X�X�m6��gP���k�����A�����7V��!�5{׻~����,V)���@�@�����d An�>�u��X$:����$�j���g�|�<w�;aB��/[��n�g%�UX�"�>�I������;���y���bOp����taHw��W��SW[�-�ך�(�[��h7�_��+��;$&��fF�]O��* �=�=B?ߘg�>9�r���N�`]��>�X�ae�[aX��y:��S���6;��kv���ZA�gI����]{��O��YW�#��篐o!z�dE��i,,J����c���rM����E�§9�@{1an#2?���`��z/n@���bs�2��
}d-�[^��Mgb`c_�5��Dٷ02�sN4���7��@ �k�1tT9�׋�|Kh�m��*�AS���
0u�z$�ٟ����:�n����C�O�sɰ�m�lv������ִ�Iߍ�exx��Ue��=+�n���}N���K���qh?��z��G�WqES�������(��Ҕ֍lW7�Rٴx:�Z��T�B���wUM��ߥKW�Kg[{�fZ�d�q+���O�q}ˇ����"b���'~�N������\����Uz8�V"b�fɺ�[�
�B�A3L��۷�������sޭ�y?��Oؙ(TSѥq.�i�6�s4r�>��|�3~y�u1�5 ��L�8=#���b���?��������(�$�����v�n��@���0�YH/o��^������/|`�Y]fa��̅Zt5Sӂ�����c2�	��\���&�]��n4�H2KS��@�0���N8�-��a�/ih��d�&�x��?�����{���m�#��`�\7��|u~T�S�h������#E�p3AK��k ;<�C����}����~����I�$�x ��$QĀt aɖ��>�RǓ�4}�Z�j�
�7�yPY�vu[��P���@���6�p�2O�����O'3�I�G���4aZ�*+�B���U�FB+����h^��V��z���>��K�����r�R��k�
S�Z�2����;��Q8�g�q	>�7=WGz]¾=��wa�� �|\�l�527��5��/��!R3WQ�>_�� �@�9�cV�o���;Y��i�|�?�=��~k��_1���t��6T\R9Z���n_�h,�C{��fgXi����ƣ�?���gN�L.���-+���������2��3-e�D�=�PK�����X^�3�Z֮*��������ĝ'��`���힪Y�wOY��]���.R�o���]�����'>������Pt�q��5���,�޺��đ�놷��,c��#�Vr����*��
,聉�Ͽ��x���^�H0F_�_�C�%��N������;+t2v2������n�.���<b骷?����
���D��)�`�a/�x�zE���q#��&N�Wm�vuy�������ߑ�Xw,-i��� ���a����'-u�}Բ��r�[�?ne�$m?_:���h6��O՘mP1����	v-LܻZVrh���ai�sx~>�84ݦf����>���:v�g6%	��Z ��g�P�i��o�ψ1��:���3��m��Tb�#�e���d��%#ɾ�%��o�c)c�A�!4d�FȾ�0C��{��s�>�u��z�������m�����ѵ����"&����@�z�,Z�P�4�*��FO�L@{[8���z塝��[v���f{�w,��ݟ��ܾ�S�Ö�� �'��+�1w��Zd�ѽF0�om�{ �T R�;7���&���&ںm8(چC�[�bO[=GD�Tj�Yp�rK�h
��w?��w٤��[����,Ҁ\��t�j��$���?��I.���K���OB5����yF6��&�\���L){H6c2����mMK+lO}*s�8w�WPvv"vֈ�#���Ü:�����݀3�<YA>�y[��[��[=�S:߉�OZ�0kh��&�9��9�.;Z=p|�MJ�'����s)�����	2�l�e���f��wR�c����X}}z�_K gG��C�WY����N��Xc���r�j*�`���i��^��YJW��i���u��1���K�6�������\3󲶻m�5;��Q��&�'� m�ЃK�>���SV��MN����״T�1P�Ƣrrȋ%G�4U��i�J�Y���M�~�������*�G�^���þ���a�f�o�#��N��M����)��j9���i�+(�H�ެ�?��(8v���g�l���b&?���-,1��%�C%��7^�.�$A�3% ���z��:wGQ�놻�W�!�4��JS.������-�t�����9���G�����E��$};�_��X7��y��6#R`��J{��v&���'(��ֳ2C�W'r�N(aK�-Ǜ.���ݞԀ�������μ�FG}ΰ�����&�I��bc��Ã�ߦ��x�������7֙��ź���M��:�t�o����T� +۟Y�(�x�{H�?������Ĭ�9�U����wP�Q�c�+������E� ��fj�����(qQ��J�{q߱�	=f��*�,Ŧ�X�����}S�6�H�	Q�SBC�B_�s�+lW38|.3+��C�998��T�<=C�YR�9r0�e_j'222�<��r�j��ȯ{���🲪��S����<�ɦe��ջ����7=6~g��.�jK�[f�����H#�����(��	��%���@ߜ<����|t
���{$�{ݺ'�`S�/�/G�|d��q\�^����6�|J
-����]�������i��5�c�MܥH��0kaz!��ϮU2
���Ss�m��q��޾��J�"]��U��(a�б�xe��'��^�r�5"b'�#�`�B�g][N7<Z|�	��b�h�b� ��W�f���n�|1�yW��q_�[m��t�J|����}�KEΦ�[��2څy�a������=J�H�v��wy+Ksw�p��p'�����/���_F�w����<������џ۴&~�vd���R!��ԉ~����ػ����f�k�_�<{q�Yc�{�t¢by�+D���>2$�T���M��S��\}�/��kym�ڋ;���^��<�"�:��^�������H�t�J����ջ�T�ޝ��G$P�@c�|U��# =*炟f1�M>���ap^c04�0N�f)��c��(	>�/�{�-j�Y�Z_�x��_�R�,�-&�G��0�#,2�Yț
`���5#����k�7'W��{�uk�z9�R{v���'*ZԾ���*�ȝe�~�0���w�{�?WѬ���xX��G}��ڄBu\�g��)Ȣ�h�S��OB��N�a��5S
�թ�C�J,���6�哃���5: nX)pkk9�j�0�`���ưp�d�d��6��&�8_��~xߚ@����jA�/M~n������>�b�9�êt~Q�J�'`��=�Ң۸
7��>�w��Q�TɄ�ӕ����`��4]�W�S'_`)dҭv�C�Hָw���I�$���fjw�`�ߚw���n�fBWt��Q��{����H{�~������O�`nN�Nb@L�^��J��1����M���d����~}��"�d��86AE)�j.����&��L�ڴo��uN�˝�+�v:%&�4��t��L�-&��^xZ*K$ߧ����^���Xr����6�w��:.,I�Z�'n�6^��DeL� g��!Z�h/��T�G���Õ^� ��=ւ�*����5�9;?�!�uŇ�y��d%�bj�1L=�W���4��Aj�_[Yy�����O;G��u<�i�OU:�/]�Z������A�̟T�3�/IG��n�K%�6.X�Ȅ�o[����
F���oE=@7x��6�f��>��cɏB�!�~NY��IyG��N��N�DjMD'8�œ��y�~H��WK�T 1�~oR��zn�n���Y���)m�^��q[���J9��D��;j�h����X��_�����G��H3�Ʋ'���k�6�wNVk�v�����|��:�����G[=�G���5����8���vҰ��7���:�غE|R��%F���,�� �Ɇ��~�\8���� ��d�`ڪ�Q�9H�>�	����Ԫ|��Y��	q�{�r�w����H� e���5�I��}���K'ȊZ��m����pC��Z762���|Fs/���Z�h�����/�|��YQ;-��5O��aB�=({y(.��
�ʾU�r_-|��ghasɋ�>��Guiunx--A�d��\���@���r�8¥x��*MM/�hs�fѺ�e�]WQxG.w��{�y{5�8�}y�žGf��dZ>?�o[d�
\H� �R�"�1�s؝�����C�N߫ZO0����[�U\{o����Ԕ�֒9��\PA�Yq�L�"F2 ��['���/xC:��Su�f�IK�q�r���� ?�D�l.m��<}����W�/f�-�U ���lfz|�z�lu�_���{�}�n�`Áo󃹏T�|x39ӎ-����P��57W)�EY�5Tn����ݼ�p��:>�6��Q!\V��]M�����=�>F;�Жֽ�����珯��,��H��ȼ�J���FZ���֒�592���	&#���~oߞ�l]��p��8?9*�bǉ�JOȖK����l��_�D޳S�����M4���ˬ*��kl}���6UN����E5�<��m�է|;d���,(Z�~�#��$�`tA!x��R����q�'A,Ϣ̋'�*d*s!�l���]n#��0�M���Cbcc���B^���JF�OK/,�	@er_h�xH�W86�������d,esg�f��x�Ʊ䣹�k]��S�����V�u��!a�H������b�\�?����st���?���F��Êz��5�/x�$���AB�]ʵ��W�l�f���nǼ��:��A)�L5��܍��8���"���f3W��c�	�����Ī�ջ5���aٰ�8>`�;G}��cq�XA�CMPxpY]��#�l/��֖�T�	�|M�t��X�tZ鈫v����;(��rݙ!��4��3jz��/h.��h�;Y3?�~�T���o��i?��=�<�Z�2�D�i!n�ܥ��-��{H��ka`�}mڽ��~U⹑�\ ��v0X◼ޱbP���t�iIL�wOq��t�(�S�H��o��u�3�.Tw��PX�u�hC����v����g����R�r����dt��x��lY��>[�����ԝ��t1N�sQ(!��ȏH$��
;�l&z��q4� �o9��A1)��o�-�)�ϡ�G���A^��������"����oY"��-gL[����i�*d��ǻ�p>J3��F�w/�����x߻�vL�K�<�SU2��C�����<�{��>³��������9�cSR�`	m�C ��զj�ۭ撝yoW[�^�NI�UK�9��Ҡ��6���<b[�d5�h*�'�����Vb�APP�Ej'��\�5�D?�Z���8���==�g���p�� *�o�r��Ը帟���!�:�g�b1�������4|5+��#�� �fťE{���*����� ?�3�'�?d�a�"fŦ2!ٌ	NA���en������ {mU��WH��'���ȚYV}`�|�ǽ��љ���>�<!� ��7�z��9A�!��(�<�7��-�H�N��	���U�t��f�/�+�U��%c�'JB�<̿���wp�?+u�lJZ��h���ɰ9+˜ 7VC��oa��^^/��P���5� ��	M>ċ�f-a�'��)>
9���>[�u�i�"������o$�D����_~ߟƘ�*)��L%������CW¬92�ږ��>���M��as�J 5��m�=|E����@�%T����4�	�qw�����ҦF&ˈE#h�[u�PS�MӇ~�o��}�O����'�P�[M��hG�b�D��u��w5na�̵��`��9%��LZ����Rp�$�#��b]3��۷,��=N��ڍP���Ѻ&,[�A{=�%%����(�i��(�8ڽ�!������������|�h���
����־��B����ۗ������hvJ�cj����	'c.A�ŭ;b�.�w¸��3�!zô p�I/�q��gz��d��UW���5���=v#�"Ë��/9\I��~&�p�)����� s�hrr26�D�����E����2{e�Ü���sr�B��/UМEY���=�f4sv���T$�Z��E��=
9[_������wǬ6�m/v��/0z�ॸ�c��\9�
zR/�}�s��P���k�q�wC�5�`�#�2�PQ1q1hs e�o�&R�u��%���dW4�P�^?����Z&�e�q�X����t{I�i�	��a�wi���rZNz�N*O�"�O)�b�Ǉo�,W�8��r�,��\��\][P�
*/�2����A?��Dl���=n@��c&�lM�}�C?.�)aoP�߲����5:����e���Z�F4��5V��⵼��a����Q-��*��
de�'�M�?~�#JϦZ��*%+��o �/˦�0��>��+)��!8L��!.��U3�:�R��#Hi�� �F�N��a���'�2�>2;�2yd��p�5T�j��I�׮FI�mW5F��xz���J4ݸB�c���x��&�wN���*v���H#��;����7+���l�I�x'���	&X�Yl���j�w�b��1m�9��v���C�����'�]		>�q����l/�
yƹQ�:���s�&��Nu��ē6���{>z�ߎ)VO ���t323-~�˿�6�����P3z����i�0t��^4�wQioļ�1���H��{o_ĢPs���f���tr�BO��������l\1�Y��BE ��3µ�����鯦�gM]�s�?C�u-_��sM�����+�7�4I�8ꨟ�δ���p��{S=��q�&!|}zd�@r´�m��=�ٞ<_Ɇ�L���LH9��(�O��̋F����X��w���s�!��)�t�
#Àk_�\���|���ha�$,��:�IƵk�1f��H�l^M���'�>%^f���������cc[t_al5�i�ӽ=��ԯ�ɗ.���t�}���7t� p׸ÅXG������S��09s7��Ms����ĺ�ٟ0��ǌ�!���&�Og~�_+��� d���.��ė��ooo߯l�go��֝42�J�O��N2~R�>�o��c���Sx�~]X=���͝�kd��[���+��ʷ��9�MK=6S���ͭ���
��nrK�K�!q�M�z5� �Jp�ꖱq_��e�r]����y���	��������)}D.=�L�yά>Zko�2]����((j1wK�;���[p;x�����`Jb��Dy�����m��ޫ��/Q���6$_winA��B�g�!_l�q}o5�҂$>�l9rN��in����)��vZ��VC��X��B��^������v���2�~q�
N�$J���t|tt��d��B~�L*GOi�T�<���x�h��|0J�4��m�JV�n�R��V�2B�;4��-<���d��`�/�&�E��S�Ns�<���.̈́1�Q���"12y�}�zl����O�V�5��1a�0������X�&�)�@�r]|����]G"�6�9�Oזxw��k)�!V���?x��� \fzY�1x��#Z6�,�N��߉�_�d�t{���>{-�;�Hs�?&8ƚ���ȷ7(1$���v�`���������<f��L1��\��h��Ih�s���9���Q��~r`|ަt�w�����(������:����u����jڌ�'5�i͒W�g�B�i�aG.X��Ġt"�"���J�^���Rg��=�NK>=_=�t�>n�i�Q��=Y\�E8A��y��+*)%"�B�t��D��'6qf��F}~��+JP;�5���gHp�2�3z!���V��FF^�_9Ы�cI�^݁p�XQ�?ښWY�uD]b�	+���X(v����z�~�Y=���w�a:��A�J%����]\ @J`B�:�����������S�����Y��S��Mk�� �Fwa��Q�����n�2�?��T$^8�<�����[�J,C��,��x�̱�%i������	x]A�����M��yj��>�8�x�;e�	l���6gZt�K��l��Ƶ���F���1u�E)���h���l���[n붜%z�j����N���kp���(��Ԍ��`��g��+�����"@��������O�1�[�T��O�ހ�Hk��j�'sѠHȂ)I�����x
yҵx��I3�#/I�ŋ�����67�
��X����k�i.E~����NhXP����w�&+=z���o؜����]�p�8�)i@tp��k���'��M��|��Pzbu!��� N��Zy%��{�q���ZYAbP<�/-!k��ˊ���
�D^��v��
���~�rr���$=�0T*{��עwx�e�����W�y�p�}|}��p��[ː6駋���V��?������YV�_F��$���K��%�O�V]�qE	�f4D`�޽��k���o7��>*���4#�?���8a�8i��P�p�~�wB�qXo__��g���%y�������`����f%�Ѻ��Fb�V�%ף�������d2��QP��y� ��⿧��V(��-�Ʃ���𣒈`Gǹ�5����qP�E\��Sƍ�
���t(�0r�S�P�|�k0ty���C�hӹ�nZ`�2u=�Z���O�y�5v�^�������f�}�[�NӴ�'ډPF�ˀgڲd�6����K �����.Sl"�� �{��jH������'��*����E]HN1H�g����B�۬8Y������	�l���rz��,v2��Ǻ	h}���:]3�%*'A��Ѳ]NGS���9��t �MB����١�����vw�%M�&�Zv?Z�-[��+�-F����v�+�Jv�֙�5�����:�K�$8=M&��A�2wh!�%�0�<ꥋ@j��܍����j&n��TqEkP�f�ۊ4FP�h�8_�O*�� _�9P@fe�nx��g����@�x�ϟ��Q�J[m��B�?$��_�st�P^�p�_��ܯy��j<��&�W�������?��<45��6,�3�r��Is��{����AF��\�!���M�7� �&$YV���h��?o��9y�]�luno�>��I7��ς�M�Ǜ�q�JVD�P���5��W;4\-����C� n�~�`��l����v���.��U� <9���ebS�ĕAG�������L��h��A*�ڑސ<{-�_���'-3���{/^����8D�y�n-�Aǽ.�mĬ�s8Jl��\l9� y���r_4�j!�U/��.&JG�	��i�S(b�fSfh4�<��-S��bܤ����࿖�BLy!�>\��D�܆�Kay���b��;`���J��"Y������G�n�ƵY?��ˤhA <~�3�������Ih�KNN&N�p���r�m��A����i3��������]�(�\�@�X-��E�S��o/1���{�[��?�B����<<��9u&뢰 iNzNB��ǟ�*��"I�lt)��	��t�O�PR=z�P�N�;/�L,��#%.��qI��mM.�>��RXxk �e�CŴ����v@[����ٛ���Qӎ�TVJ?����:ML9�܁j{NOWTıy@�P5���}����n�y�k�aڗ���P]���Qh�}LT��(�tlc��̽^X 7%��q��y�92�,&M҃<HMYz%~����W,/���7ﭸJ@W� ������{Euሪ�j
�7�WC���bW}�|�(���kxQXQՄ��M����;j�߉�>��.��v.m*v��2��LQ���@�:�C�P�W3��b-�����puO���m�T_��2I�/7�hu�5L�M:�OW��kqw��#X���M<�����陚�Z���P������d�۝_�ȑ�����o m�>P��g��!7D8�T�\Ðpr�l�r������DG�	Y��Ho�I?C���t�r�����ƅ��^�w f�ǁB�]�M~�]FT�;��i@
1W w!��K?�܀|��0�u..��:l�Ⅶ@�Fh[�s*�	�L�'�Fʄ���} ΄Η�FF���{�H��ބhPMSS��̎Sk�?��L�����b��u@����z;�w]tSo�����b�b7|��������L��-,cPQ��:��<ܗM�QV(-�n�SuF~5m�`��ɺp<��'�D|A����r≾DEAg�~y7�|'T�(�䵃A�G-�&wx��N�XXxw ��Wq���܈#��O|�j��8x��=K�ڨ�y�Ȉ��r� �K!ʫ��:��ZBB��olP�M�bbi�6����*ѵ�����ǩ��������œ-U⌵��jf�J�
��G���!�N�[��$�I��1�@��	�Չ�m��Yw�h��a�u�K=p����{��Wn6�ÓO?p;��PPiz���T�@*���Ǐ��� x\RG�ƥ^��O�L���	i.��c,<W��m�?ũgݺ�6�PDAg�ˆ�+B����}*��|Z����a�ߔ03�,6��mG-]K�(O �7�I�PgJfl�}�`Ħ>l�+{��ܺ���
D`�c���x*c��qy(?�bYه'�+���)�Ph�2����:
�:�huv/z	]�Q �)�5�5,�3p*��G,(�̘��$���]�:���D\G�ϣi�5�@�V���H�Ry����N��<���L�_�ě��������߉�y��6l��u��⼩�4�;dW�<�/*����yq)[b7L{ ����S7�`�p�/��x����RJ����s�rk�{!��j.zq|�>���QXYY'��@ƄV��+hk��f����ϺG���ՊL���@u�����Ts�K�6��9��r6�%n+G���\����0��W0*H���o���5,� �y�x�}+6�6U�LP�<3`�7���}9�B<��H�_����)׀f�(�@[���*�;(�s=�Ȃa�W�k�ĵ��F�_�8񺍨rU��"������Pq�c�C�ϥ�B�ߺtG����C�W��	�+����ݍU��Q5� A�9��%���
~ePQQ!e�ɀݬjo��Ç��L���_��{m�ޯ|�V<Y9- �91�&��A� �{�!���柈BhBł�����Z�

fzW��Z�|�`bTo���'�3u+�00�3�5O��v�xD���j��騋������Q ���	��
"4�4')�3�0_4�un�9OK�U�K�۩���sμlp�m
���Pc"�a1��3��.N^���q���	2��Kg�D�C�t�K�e�?r���ݽ��%�:Rh���~��.6q���zL�e��'��a��Im�I���ǧc��ܶ\���tP�v�?Ը�h}��!���߼�,����ش��:�N�����ȸ�!�uI�ձ���+D��/R &GF~[I���7X�M�]�XM�� ��y:?Q����bꪯ�Gu���d���>g��l��}�@���m��7p-da���{Nyv���Ƌ�*�\FY�Zٙ�a���0�뢑��x�7i��Cq�f�iVE���nD�{1$�u"s�ِ��������@�_�^�;��*@u��q�xtܳ���|�_.��T$��B�K��-��5��:N�>Ò9H�Қ��d��A٨k3�2/EY���}w�-�[-ٜi�ȃ��>�n�m����H<�`��Q8'PZ&�%>�U�zԳ;���}��۠�@�E�	�Еy��dJ�
�P�$���i���st2�~`��[���*ɹ��-((h6�,㢴O�$��T���c��|ZF�����28B����L��&!a���n�|I�|/���fSA�"����n2������U��a��Ёu����5�؎6_9��(�ȏ�k���J���n's�2A�w���4	�Fs`a���|�d\�m'd'g$�Vy���<���^?�ƔFK��N�6Mo"W���&�^M�M?��/8�W6n`d����SW�!��>;S̟uS6g�=-ܡ��'Q�G绍J���J'g\b,O���y*�1�8�~���G�5T�tD�Q_)��[�{WM��ei��q����Wy�	튊+���\�����L\+j�jO�7=�K/^����IMP�U�TnR��1'�m<Dfp��6��ƃ�͹�V�+�a	΋]ļw�Q����O�~r���1E���.[?oo�h��	��|hhh�"B[���L���~�w�GL�����ܺ?�A�1�A<Ln=�:�1�z£;��j��!8�! ���W��D��(����q��LĩC�`��>�~@�5�}��w=,.��tfTR���	���(�I��\�:�0��y�j�R;����:�����w���!�!�����as8�j�_	��V��Lk���[�3})��'7�V�|M��$v��.L�a���cbr\}*���L9j���**�+�s�+�L�k�6o��x8�S۬w��	���n��򄝄drN��������MzaD�9ұb�D��^؍�+?���ptk���G)������ľ�թ4J��\_�<!��o�
{��}�H���3��^�F���u��g%번�ǻg8��|�R8��~,�l-�v.����!##�����v��M;}�F���P4�6� �]2�od��9b<�V5��j8%,6Y.��Xe�:�7���OT���z|���է�Z��o��̈́o���� y�'�ja�i������}pBV�N�dB��F�Ʀ�y��)v��Ik�7,��)��G��"�9�<�K��#?�/"�>������Iڇ3>�y��c~���U� �G��ۨ�J�D�0(��E3���s)(jQi�� ��6CB���>dIxǋN������-��ܿ!��౱�Nq�YŦ��/���nM�����;t�~�3->�5Y�V�P��ن��j����B�d���F�#�v�v��<�k=����Ϣ�2IJ�Q=��Mi�U�(~��R�&n����������49q�ZL牭��s�$�G�1z��h��P��Q��=�]�7���G��?#����,.�>8|%q%�bx|\=���3�cg � Lo�ӥ:���uB8&��ڳ��l��W����ۿMH���Fڲ֚��MӼt����
]'��aSeN�������""O�H� {�:�2�����_��t�_~��S�--d�r[N���l��wjE��N�`�������KC7���InY�Ͳ���Ж� ���q�q�ӹ󽈭��V˃_�����{�]��gQ���dc��DԖȁ{�����+`�J\�~Lz:"y�6;o�����������ek�'5*��zH�mt�p\ ~���]?��e�l����G;����I>�:��Q ��h���NVX�Nb�W��YL��.��{~�ֵ�ϭ���6nݛ�UU��)BՓ%%ĝrtܟ�&* N�kg��7!�B��Q�O3Y)�r�f��5Cy�I��T�����P�;�=�5�#K9��{Gv9c��S�Y��,���n�3���켈����ϊVsJru?�����#[��)s���l7���	�}R$	nyP��(Ϋ 1�ԕ�ăKQ�(�|!o�ɏ�qB+��[���T�b|6�
�Cqi�㹀�:L�֡�F�v�\�#�*�Tk��E�c��R�	;���QK��yά>2��MD�aF�P���Ү��� 2A�/y�F��`��c�A;JF�������{ٶ�t���9!��Uf@_�9R&b��V����Y:���׫����IW���E^���"/�+�[���/��E�g;��*�L߃��	X��ვ��b���4��d�+��q������~�� 7J���oɎ5�m{���{)�nw
���߿s�Qk11��}/0�j�<Ĭ���;�PO}������U�T��&��k��;��"�fJ�!ꎞ�nu��>��؜��C��uBW$��x������c�1}��?j���㪧�(�����I�y�q�Q������}�+����@����%���t��:�>\l ��9~Xˈha�h��J+%�,s��WW؃��و�6��HDŲ=�*^���G#��g��8��+3�$���-0{��E��j�ί��jQ���4YK��9ʶ���oVq�|��D��$���&�) ��Z����RT�I�K"He+�֍�X��������\�M�/��"��Uqi�7ހ��aL��9Ʉ����ʲ놰���N~=[��_R
)q�D�zI��~�vp9)�n�����ֳ��,F9��ڻvd��7����2S���9S�$�^!���D�����n�,�	�f2�[��-�7.�/�X�Q;,��$; ����c���P��5�a �x4d�y#�&�x�@��:��eV)&�{Ђ:��v��0t�������߾([���7���<�k ��WVz�=Z�.�kKz���z?D2���[��r좗��E:�5r��U���Q�ޟ����U���̧�r��ˀ�a__����*�T�).����	j�ʿ�����%~���;Oa�=�K������N$�X�geu����F���f�%��f��K������W)o�#r.�.v	%�ѷ�{�#yĽ�H}��F�e_)��Qa�G��0��t�;݊�1I��k?L�%88U��
%��9�����FU�֚��ݼ�*^�����A�*�7�~t�����٩ ����K�� ��!l/t��gQ�fl�[�0OVL���{ '��4~���Ǽ)y�7$�<
�p�)'�I5�4|�4��w��B<�$O���\w)vȲ��Z��B�_�M1 �u�贯E�
���[K���N��Go^I|���E�˕���}<��Oߵ�7���B��~��_�����ي�y����Ӥ��۵3{~�2��l���Vq�ǍM���Wo�5��o�)	;>o&���P>l�G� 
����;�'f%�:�$�k�#�'�ْ�Mް��[�!2�Sx�e����~sG�5�ۙ�kqѶ���&��-��(����̴���+̦h�\�ᵂ��B(�Zъ����~Yb�~jї�L�	]`f��B�!7�}��g\���T�X�q�'�v�ӎ%rgB�`#	����W4�.}�qy��Z����UTP�.�Z�\�4(3�]G��2�D�* �77�ا
�f�7y��ǝ�ܳ$�y�F�P��+�B6:��:��E�/��2��"�%^���h�ʄl�*�|i��(|U�{<���qI�|�����:(�XX7�?v������	���/�m���R]V33���;�:�/��L ��(��>Q!�L�ʃ�r�����T���^M��5��1�I/��pz1:����'��Y���C7*̟��ٗ7vU���5K3@
V��H�hR��=��n�5���!�Sh�P�`!1/¿I�9�/��Y�{���$�2b��
��:�y��v�N�����qy�����	�*@����ˠ-f�^�b�8E&�i�<��.@*|�
���6��ɭy��#0מMe�W�B��8�(��a ���o��+����{����Ul��yCC}���Aliv�p�鎖�ܸ�C�5��w�Υ��μ4�qn���2AF�pV	/Fjf��S�_T��v����S{���Ϙ?�h�\��`iFz�'N���_�_ݬ��۳�x�,��%��D������U�I+Ό{�ka5���ҝ}�������w�ws��#/y���F��#���I8錎A�B ���F�9! 3�����RF��(�3�ͿzHR���B�/kSbx����\�
�N�#�	KU����r�εh �I��b���.kIB��/yi=M��\�p���z�FC��xO3?` �&#`w��   ���c�BuA1�Y������tz27����uɤ]�)5`�&���g�9O�f&�H�)�b�z������T_c��3Z���#�4����@���оUXW5̕5�l�I�h`dԷl+y��:��u_�
К�ύ�;�/�Ӥ��C�*�]��S�m�\X���)��ȑ��h�c�NFFN�7\8�M�����]6�He�#���O�^�O�vO�2��{j"h�{�MW7����r�-�j�'�GA*wCHaH��o�u0���(D´ҝ0w'�n�r}�~9�S��qz:l�`��DU�n�!��dTb���9��K훅k ��GV���, 3>J�WO~�u����v!^�ĳT+��0�#Q�kX���(�x;���.�	��s/Z���ߡ����sy��W��0�WA�P=�d_�x�N��`�6���W-�f.dĭ�[[ie3\�>�}����I�Z�H���3���n�Pܿ��z4�~���ݭQ����h�m;<�+!�쑰^ٸ��j(4+����u_�m�WEkkRI�D�9
ІH���2����knt��a�yEw-� ^D�2���v�����+Q��dr���m�r���%_��fd�6G�������w�i��-\��d�z'Y��H�����H�F�cLh!�v��4�"\Ӏ�Z(�M&�dtu|�׷���:�� �EYQ���{I��hʋ�qo`
t�bQy"�dB~kMU��Ym*ZRh �~�s�)�/hr��˻k۸�@���I�K��U� O?���Y>����<���}?؛�g�k���Uw�( ����:�ܶ��0�?��r��m������֚9mv��* &�ݤ?"�)��j������\
��6��{��� ���܏93\��7��Cz�p���qd�u��}v�����Ô�@�3���?��q	P<�5�����+c�����c������	�]���@ �Y3��3�~�E_"hu֑������H)!���W}�^��Ǻ���s�P���ha	���͉w�W17w�sh�ы2���B�(��ywg�R�Ix7"�'Q:��x=�H�)l�C��N%�)�,%����5i��;c�G?ŧ��TǙ�mllL8�==����ʲ�F#~�/����������> �h�)?3}
�H4�L����\�����N�oD
���o���61s���7��?	�ϯ�a��(K"����f�QCkCF��!��sjj*���/��U����
��7��mS�{ՙ߱Ӕ�M������B�&���	!������ڐ2��X�3s��@��C��ȑ���J����ۯ�$Z����T�Y�����Օv�+���暞�M�ɇ=ΧS74�u1u�f���i����T���
~���S=��U_0	��F7�T�E6 �9F? ��H���[��5*��zL�6�M��X����S��핅�
C*C�'x_�nA`����&� �
!��Q����ҳa&�����A(�����}���|��(�{�y�{��gdd$t�J�1e��^x0�0A񽗑���]��ώ��Ĉ��{b_�4��g��|�aS��bO���SV:�����_�&�nE��VUL�#�̼p߹rm�b�qXc'�M��Up �O�:�FQ�yA'��-��$e��\����O�WP�W��W�k�?��<��7��SbJls��B)&1G��#�}_9f�[�Xs�9C(�#7ab�\�]-���������y>����|��籶v�����/��FxE�b@$)�Y�.l�}�ܐ�b��W��i�"q�J'K۾��Ƀun�W�I��ɐEU�F�xďQݙ�3�Pq��-q��SB >#�)���r��
�T� ���ݟnx9E���}qҦ�L��K���I3�� .����-���u�Z�$���j���-���º��g�'�U�d#)��`j���R[���_\u^�8ɗ��@�R'?���S1�J�]��+*��p|�A��a�յx�Q�ʯ1$.U��& ��?����{��LMp��[b�#�XC��@QQo�Ay{SC���TI#�ﳆ���?Wve��&��h��^;�frb���ߩl*�&h�w�>r[�I�H�}v	a�t����Ӎ��R��w�"�S�mqQ�X*�^��[Ѭ?�f������^=�'x��s\���(��}��jS��8�R�%�6���iW�^/��\�^t�_,�^�c�߭G��V��/�b$�N ��.���Y?�	�󘪻��^;�����G��~�Er�0o5�,�3���*%�(v���v�sM���Z���^=�Z�?����0�>W]��g[��6Ҿ����Γ-���������T蒾�o�_~N����6�\����m�����aar��G�D���o�jߴ�֬f���X�i��i����MY���v{��.s6�S-���&�w�lҶ�l߱��oD� ;�G����]~{��@��ty�ߩ*fE�Wѭ���C�T����w4~2i���l���s^d.�����h$�@�&���b���]����B�\	�s�)�q�6��7/zKT�H�t�B�ϱ>�jerE^��������V��9���W�v�d� ��J��<wJj?b77�|��C\OJO#�4lrlƌ�=�� 	��sW��[�'H ^�0n8�
?���綶J=�j��ʶ�N3,RI)���5?�Q�7��)�wChMd�+�`�HE>(��8W���Qq�Ra��rI󰲲~Y,5z�i�9ܔ]��3YR�u�����0N��o?��;���,��\��.�`i��A���ea8�
ig��2w�j��V��;�"�v�~e�VG&���h[�{����;^<�Ľd?9�آ���D,N�*��K\���D����YLN��N[g�J��5��Xx�m�ɝ�T���x��xs��	8�VK�c���M�ʘ��v�n�鐒���u�]��?�~�ޱ�1K���aa=�o?&�sb��� ��Ģ�GTO��C���SVZA8
�	���0���쵵X����zZks�Ħ����H��?���7��M�??��K<H6u �A�\��%(�(x �P����x�)rv�\���� #.����W^�ځ��@ �G՝��"��c�!��e1�KP¢���|��mm9Z��h�Y�q�d6F^v�p�l�W����|�?���K^	<�������ֶ��6�����Xn۷Z��r��	)Ĭ�1�ֈ��0Is�R��ch�v�v�X�X���m����fkF���z����E:Zf䫪�a���tEYn�>kN(�{t$�5�0�\�l&���\(x�؟0�z&��5�F_�M�l��D�):�њj*b�晨���^S嘡+N����`l��B!6����عIk�ș�PjcF��l��}5�J���>��N?9�;��`�����lNgЗ�r�T��������kc��V��'�ka�ӭ�orU:�U:L�:���v�1�7O�-��|�w�����ǽv�i���Ѿ��U�1�$JK������	U����+��n���ߺ\�e|M������ԓ��vs�ڀ[#=�h�5�f-�m��8����rވGx�ҕ�� _��K�b]��@Z�K��
����I����O�/��0*j92�Zp�P�\U�;$�z����^�V(r#�]�����v�C�\NI����m��0�K @�A���?g��?�@@
�p�΍�1��>�cZ���՝��U����c��M����?�����멚Im�3ָ?�qɝ�\�GIo�NQ6_��M,G���=,�f�������gim���n�,?b���ǲَ>���6�X���%K�R�YݢH%�	DM-�,{�g�̮FG�O��v�P.��ϕ�臼��F��`�.od6�v�^���v�A�
Ϋ/�}`+�k�=�T�6G����xfk8~5W��X H�%���c� jY��E(+�K������ڞD��} ���շ������h�޺�$A���0<*���z�|A�6�J ��_ig�W��Q�b�6@Yk��O�{$�|����oǓ���X��n���z7�[����/�����j#7�Nc��F<d�GB�����ZvIqL�O�Y��o���U��J���JZ���_�:�*.R�W�ڬ�ȋ~��F�)�NXv��k�÷�}.�`���%pa�~ TԾX]�]��%K':<r�Z~��t�f
k��/���s��L��W�:N�\�y=f���H��됇\4��y��Ƕ��T[I�冿g����֊�e���J�.�X�I��}u>�}�N�K��1w]���e _t��m�,��ܘ9 7�Së>R:m?57��/~�*��ۋ��k��2��P�ʳ�͒�O���n
P������7���8��$�<x�o��%����lf<4���ϫ ��ܬ�_������
1�w��l���%�+)7�\���<��AW���!VSު����9��c>���P�l=���m"��z+�5�p�|Mu�b�$���"@.N��`�~�eX��)e�y���FZ�P32h>����m��N��3�)��']�Nl�ݲ	�W��	�������kC�~Q/kn*Z�5K�gڔ``"�|̩�B�ꁯ��x�������͕]X9g�z(:::~��I�۴�6s�Z2��B��6��bQ7����$2�"9E���]M{�s?WO�Z�<P�����0��fyy�����p�2�_;�jo�ph�N?�R:�a�S�����	h���h��]�;'q���J�ӬĒ�Ņ�$�;�d�m����F�\��e���rKY�k
{�%O��2�m5	�Ve��^E�a9���a��ǣXs������ZKhxxq��\���03�W،��+�N�75H�$�I��R�?��/���II��7�����;�ts���W��ȖZ)AkD�t���6ڹp�/н|����[D��9=4nıy��K�``�\� �p�����۹|�����8`*��P�����S_??��K�fQ�b��!G�b�:�EW3@qC�W� �ak�2v�!��}5����9������%���P;�ؗ���a��
rA��v��/r�)�<K+���e�Pt$^�����R
\���?v�~ �1�o���諱Ǜ��y� mvnU�9 ��߾Zw�"��t+�&�#&���"/�_�آ��c�6�N��`|q_���#^�l�o��M����0+�����J2S������}>���B
�����n`Q��$f��8��#`��ݦw����T��M�ͰE=�:煷>s�"q�b�d9do���8��p0�΅b�c|=p�፦&�����J�ڷ�z�\�?�j���}�r��*�c�ᡙ�"ee#�}�O6�X

�Mw�*�#��r�$P��R+��KţA�#"�ִ:�ྐ�g+�J7��Gy��.�3-w��[PX�*@s��S���Ô�Ő]��!A��<����p��|{{D�WH-��*Ԩ2������<�;�Ϊ2��m�j�����"�`d�����<���p
m-�X���pC�s.�o�s4��m�pOQ�^^�[85�\�y���hr��|.>B�f���n���k�e�!S���c����e23Ϸ��jj�o+(��%s#���U Ԗ�)��>v��
o#��R���l�nh�N�.�#��ɗR���}�n9g޿�9��~��o9�����v�	K�N4�*� ۏw��*9���Q�R�V��܄ }^����ɷ�������5������:� �?�m�K� �����-@�أ���;��0�yܣT����8��V�L�Zn-���m�iw��_����rT�C�P�-/z��)0�l���|��O��N\�o�'�K�ȕ�+������$	�܄u�$�*<X����-ڳ֏4s�����˚\���	U�������(�he;)T<؈){k�U��=׾s�/��q�,�G�6�����asԈ*�����V�=��G����E���WߣKVZs.i#z2����Ĉ���ݵ�-���37�a�Y+�F㕨ݷ�C�B�1����\F��>������}�<��Ԇ���$�~�PL�s�%�� ƥ���VVVޤ-V��q�H��	BT�y+��Gq�s�4ƥ�!i����-�/@Nۢ�8 L\��d�Jb�Yq��.i�?����|4�	�<]�9�\�؊��Ed�� 5.ƆRN7�y�5��[���2���/��j�px��v�ȵY��K���[ka�����r�D�e��2� o�L�	�g���!�ZR��@�nX��G*��-:qa�g}���ZK�1�3��$�t/s�V����N�M��xͰ9R7���Ej�U4����@nȂ���$(ʙ`��w�� 3��s��l�����r�BNV��?o�� �y԰go{j��7��ZV�7G�����+i�!͸��é������3���V�3 �bg��9�{V���dȡ�0W��w"9���y���U\�^"X�=�L�ňN#�ѕ'��wI�Od�v:����.��PLu4��i��(�=pc�a2k��|,�m�wx�[��J� ��b�����6�/�N�%���8�ˁ���|m[����R��bv��4y�f+�_�#M��)M��d�Ü3az�T��춈9�۫��a�j�o�7�)=� ͳesgdV�����Z��Yk�]l;�nn5tC��r��6K�>��5���/:R�	�f)���� jRRg|9E&K������Y��v|d�E6�G�"�7~[9K�;.I-�N�C�ZRt]l��)j�W����-b9/�:�MS�\=Z�G6[�����<)J�û����P��W$A4O����L/d�4_G����,�F\�v[�7x؍���"/Apm������Rye%@�/�K0_��<a�����FYL\�����
_�9��2�=/�9�h�ܲ|��0�]�;�}�op��օ$�橶,F���붅X:��xi)�w�����g��X�Y}�şΘ[���Um}4�0�v��G5� �?��ڀ�~���d��0`��W4z:"���v�gAe��B�ͧ>{�^闥�`w-�ܫ_�9t��P�ҵ�ٍg�Xz.�dm�\�ҙSS��,ՀW�LPcĀ]}:K�VS=����;�7G� �^yT�p��Xi���d����av��#��_b2��/أځwJ}%F2ξ�zR�Sx�<�d���Ǜ�h�#"��}��`�x}���Y�܉,P4H�L�Ӈ����h��� iA&�\�v�%$��Q�b�Ԓ�g2d��%�H�\p�[5Ͱ6w#�_�����?{*��"E��t/&nM��}�W�T	�I�DjF���sC����G�[ �7KdEP���s��n~���ዼJ�r�x�yjcN����[��
�B�L8o=_'XxZ�������(7�}�3qUBP_^|%Q��W�Z��&Q���Pj�tH�����mgv7~dk�m%�'��[k�'��Y��\�߄f ���ᘠ�]�� C�r�D�s�7�?\��}x_���� L�ڨ0x6�����쿃�����V6�6uk��iL
v'��(z�gp�M6Ӭ�����Zc y;XTU!B�#��Ծ,��)�-�ܥ�,j`��F���O˴m$$��������a��6ǔ��[�)�t� w/D>��{צ���V�?��Ĉ5�jݑ�<�����mҊER�B�����rz��إb��0�wl���oQh���Go���� ��&8	�Z�7ʞm�ь��3M��x���K��ˏN甞[�_�l�:,Y�������wIB��	�Vy���.�����wH�ংg�4嚧4�Ap4U�< �����iً��Tk���މ{q� ����j9S����=���S�����go���>�e[m�T���+T.�����Cdz(��e>>p|�;"e'u�?x��.��^��\W_�_�����wh��BUGd.7�l����j|���o/�[E�wV�w u�6Z%��!�g���r�UihW�^Ӛ�O�� ��p�G@3�8�bZ�"��m�f�n�ѓ,4A��pU1B+#���O�I�~% �A�\��9Z�i3W,�x���Bm�\;�� �+~i��uR*��r{�1���Է�t���ƽ�M�W��z<Rg��\1��8n��fb=!u��9��Z��*uGi�������V
ġP�/��]ə@G�t+H����
�o�n��4ʞ�F����8m,���T�tB���r*��wB�9�
[��~؊3)_�?
� �Sv��*�I.�YT�o�<����������K�Ѱ�D��]�4��C��� &]4b&#5Y�XwJ��HvsVUUA��D5��J1��_)%�q
�D���Ā�q%��;?���<Йp��Eo��M�[�:�?&eX��	N_P��9+GJ�Z��2�������|�\w�b�����O�����k�,]�tA�Q�0�9�9FV>�rH� 1cK=Hc�\GܲDާL����t�Fw�G����AŻ��j㗢�3��,�.m3�ǭ�%'�W%C?%_L��2�@�K��)�+�^![dP��͗�)(O��5�je��zѶ���,���򜸨�t?p�7��ic��	���,$d�'�����TE��(��%55�h��8�;�6�ZM`Ӊ+4ťwLX���Ǟ�˿��FK0�h ��������(/�&���U�KM���2WU���!ֈ���Ux���hU��n��k��H���y^m~�`s`��X�w��h�n`���K����~�`��e��b�� %��Fz��2g\�(���\{8�3�O�V��G��勛<"u�m�<��3(r$I!TU�X��Ȧ��Ge�I���s���s�������0#�.*���1w)������3�V-���-�
B�����������X��,�3˒�}�]��JФ9� ��Uj��Ź�K�G��C������̃��R�$0�Sknm��RK���]\u���.y��~E(zv�P�?�KeM��C�aʣ��X��4��)��Y�Ҵ�h�GY��\���OX�L�O>Mc��	_?��	���������9��|W���VG̔��J�q"��V
XU�	�mk|!���8
�*ˎ[���N�u�vI�)��n��?��ָ�X ��T��7���PCws����*G������]��t#'��ҹkh���ƷZ�k^?��V�0JS=Y%��7����	��N1���g{�Q��R��95YA��a��d�/ZE3w��R���dz�;s���A�_��S;���Y(r��睩��a���UI��	�8:7)ߞ�v�6���}$�jUk���,��5�Й)�������)IY>�!m��(v&��>Y���L��SQ��?s7AUxÎ"$����[�Tg�;¬Q$3ď�Ľ^��*�s�Mz4�[�]��u�)Cn��jX�o���/^�Ke�YU4O�@~l��F�~~x7Π�Z�Y���[�B���&��s�=
����
'�z�2�����a1g#�M��X�8\k�������E����������j�t?tJ�'���Y��tf�X�i�IA与m��Rh*��4m���%�!h7�v�+6U��q*��h�f1 ���lN��|�%|`+�6'7����}n�3�ߊ�%1l�.�����vN�`���?�i�8�����},�J6��3·�n��O��Sl�Zk���$P���V���>��s�|{i�m�6ᯣ��꿓'�3�ӏ�[�+�ͻ 9�x�ay�dP �?��9�l8��"W�3��e��E<��T�>��	��bw���n��q�����}@��'�;�� �w�C��������rpn�:�*��o� 0i7�O,y{�˰a3�E����}�rxҟL$�ƻ^�9��"��Ϗޜؽs�^����[�E�7�5b�����(�}��@��������ɉf����l�Se��{y�|�e�K��lbZ
�����s/�e��I�t�a1�Pz�w���Ҙn�U��_���4�.�����,�����E��צ�����S� �@�_������`Q����m7	�n�س�@��&�����{�l�յ�v
J��G!�Y5�/оo�D�OF�P���^6q]1 ����ً:5�l¶��"g�� �A5G�2/�~p�� ��`���W���OFr�����f��\=��p�k�(��ޤ������\V���ʱYʤo��p�.�Gl�[Go��ޥZ��[��U�5��y,��Ղ̂��bż%ss�􋭡��z���% 0�����m��P�>MGR���Ns|g��9!|��վ�,���9u�?�9<�7~�@!��B���5�XM�u�[�"�,���KPz���t���f�a���  �j�$�(I�g�.C?�1�mκW��qPj��<&=-�� ĭ�+b?9	{��������я 6@����>Q�������4U.����b.rܬ1��O}����}��$�u�G.7
�9.8�]w�Q*�l�-��G`og�Y �Di8�M"5+"�qil[+�AD�q7֊�����%�wǐ�y�UE�������_C1ޟV�HL7�f�i��˯F��J�������?��~���rކ�ޚ�P��ޅ�?_eJ��`<�?$ �O#�X=Q����`0>�˺�z:��ۉnY��p�x Q��g-���W�����	��i�����_�k�+u��l��b�A��L{N��E���,F�� �z�����\�C̠jS���C�N,naoy����{3)��I��-_,��x�Q��C'ة��K�^��+YO����ϛ"�Er��9Y���+�6�����Cբ$L&���M�ؠ�"z�V�Zy%/w�|����[�=ZÌ-��f����`D	���]UUP�����|��p�{r���c�������TW�C�k��}f�����<�13C�g��W�{�'�ռ�+�����?���;���n$.[�Zk1vSx+ �G^s͝�[)���?���W���>�j�?�$J;��]q�%>D��_��H�(M�[u�������)���!�m+��Qq�+�G��tl�rޟg3c��N	�L���0�x��Pl�.H�_dS��=���9<�����*���^�]֝T��m☤�Ȑ���A~��������+���w�8�?AO��E��EU�97��w�)JP���{�~�[��E ߏ�Co��8ygQ��I�C�7R�.꼍��s�|�w����y��Fi;�N��nۀ������hq5����2��IS��<�S�"�e�� �(����6��ҥ���z
�U��M��U%�g��;Y�ʃ�}�^���֮���h�	���)������C3qIB8���u�zTV�R6��9.���M��TB ��V
�lɨJ$�E�o-,�$lFS�E�*�"�,9)�l�D B�(� �~�AVIfJ��y���چ�G ��>�ätXN�E�	 �u����"�[9�K���D��$ou����U��1o�_T"�H\��Wɾ,p�o�"�+�;t]��8Lk��#"}�~������dv��t �x"�s�C6��#Z��B�k��ޞ�KrL4���IQ��?6y�O.�i\�H�X�+~� �9SG���a���K������{�9����`�a��~�υ��-�׼����Ԕ&�ֲ;�����VL�v��v�5���Y�ѕ��B��
'�R�<�
j���X|�A!R�!�;Z��o���#��ͤ���m�}klr�䳲��/��� ���4��j�k�
)d��V��td�jL����Y��.*?ds�/>iq{��u�th�;��H�a)������v�������݌9�h"�&�Ϙ<#H��c�>�P1N�j|d㳫�/��F�W��ւ�)��)�y4�!BF�=���`��}3�0�t-��~J����vS}1�$�`�e��~�BY�/0F�t�(�{�d��R�9(i
l���:�4}O~�s�#XT����`��4����'����[	L����[TK�Q�5��w����{4"����V��I��
E8ʯ>����J�R���<�z_nքԚc[�l!͕&�g��n|zlrQyT�v.��7	���j�GqĿ�=˃v�%Ж���;	C�9]#�ܭ�wr(��srfdh�Zj&�M��u:��EU����\��΍Զ5�.�cD� =u�V�;�\POn���*q/D�	����~Žoe9�ŀV[�Y� :�𡙭.�.Q�k�H"�<�|Y"O��ո-�/������J����<A�67����h+���k����~�C��<�S�(���-s^
e�gF�  լ�'o&, ����>��e�ݓ0/�A�#E��[���A������:��R�����7(ha4b-
�͜���h�Nk���ad�*<�!T��З�!����G[�ޏ�d?C��go_Z��n�|8��_A���Ł�S}j�0���SL�E߄k
���*�_��#��!x��III���:72��,ǌ�P)��B���#$R"6��N1&���h&�zV<�OO�Y��W�.+��Ŋ:tI��w9� .w�Jn�sd�o�T:�N<��Xvӯ�h�G(?��um3���'�G9l_FFeǥ�?�� n䔰�y�մ�A�\@�������,L��LT�%��y6��Ҭ����e�|H�\ �~k�"JeZlyI�YA/E� ย���v�u�$os4\�"���t�8*j�8�������=Z5f��vs�P ���������bi�C����Z�L�ڏW<�d/.��y�?o<�vɹ��{���|��M7gg���ߠ��wͅ�(���y{o���Z	Xi���A�bWj^#�~EvAC�M�x�\���SV�E��j¹�I34�E\�`DK|�#lA��b�R"�Z�#p+��q{��vG\<=��I�����4E�b�5������S�`J R*oH�c��E��j��&k)  �U���|�d�x��V�sc�����~���M^ؘ�~2>�:�5�"��Hiw��x�v\���;����so��jh�QNw����E%4�jW���/j4�U����R�pzr�0x6�>�7������׀P���ti/�v�K��6Yhi��hwkG86��uf>�N�5�(��Φ#���G��ۧ���Yf�K�;@�+ʖ�����t(u��&��u+�#���[Z[Z��Ց1���dx�YU�c�:88�f�5�z$9��t�Xr:��	>>�9��K�l�6�@��U�_��O��w)6��r��PȌG�Ajjjo�?j%!^p�NWL�h/
�&Q�r�~-mN�NM߈΁?�������3��YX�E�]E��P?I^�+��v/]��Y��ҝB�,�t��8䴄O�&A8�bm�RYj��w1A�,U������+Y'1����3ml��711�jA��Q��v������\���C悇ڍ�dZ\���|����-a�N�U�!��7����	��h����"fr7�7�k.��l��a^\�J�1�`�K@�����ѹ��#��Y��a�,޶>� R^�!��@�!/Cy�{\n`�ė�ڼ��Q��^r�����No�� {�����O:LZ�8��?��_��b�t3�Nl�ı����~��$�C����� �q%#���2�3ָ��9Ы.(�S%R����|ȫC6P\�d�����H��û.����Z݃���("/A�+����X�3޻@�2;�1F�����ΐäb7}EP.��&/�+T����rî'�Ϋ-��u,��Բ��M5HC�'�M jj��C�M�D~o~Uڬ�(���!<�?8�p����{�m% ��Zڋ~���N���}sz���0,�P�*%@�;a-�S�]
Z�G �|PG٦<��x�q$��2]����Y^����sS�^�Ǌ|�c���xy`���v�۾E;��a<���Q�H��?�c5bĈC���F�>}a�����E{{{A��:�O�j�N��g�����	���褮�d�#Fȡ��������W�	�5��|z�S��ǿ�ٲ��r���^P�2����9z�k�05}r�p�ޕ���3X}(��pG�<_n^�M*�*[�s��v���M�(����8K�������ЍNJ��Z�Ν�L�X_���z�t6j|9t�f��4������ܩiT�l��H�Daj�"�rj��U��Pm�5:4�����������/f���ear�i�
] �U�o�̐j����8C��דs�_
y ��s�m��ic��~;3M�Y|��KQ/���`Է��ܯ�t؞�[�i)EC�E�ӧ��Ǐ���u��f�F�flg6X-�cQ�`�}���N���4H�5���A訞Kv� �,'�a��U�+|	% �2�g����hE����Y���C�s�FQc���#%���L���V|�-�,w�*>�٧ޏ�:S;?X�v�|�s�*v��ͽj㛃�}��w�������nM�6K��J�Lr�)婵�pWK1���
ڛ�֗{忒�Ci�BT^�W9M $A�k�
` g�����IeVm1���'.�e��+��:X__���Z3��êJ��1o}�fι�Z&�A���%(&�y�y��1�̟"e���x{DDx"��)s��������ݥ��Z��uz7�d��<���a��=���U�a�92!P�yT�
I��]��F��!omX1��9*�����x�)����X�v������V˴�_����&U����a�$��:�u�މ;�@��Ҍ�?#8 r��!�ee�t�^NaK������.mg����>�¸	Ei��)ϙ-Vl)Dl��1����c��D5�.��㔞om��J5��>��R��3{s��{�32u�jt�ǭN/+��Y������8{�Ľmzks�{a�t����,NNNڏLN%uG�Q�z��Zk\��Jӝnf���a�8Ҡ^�T�o�ӄ?�W�'�����4���q�r��du�'��X��&͉�Ѝz�l̍�YEO,�NI������Ayzicn�S&l��^�ϕ��=ˠt�$>%�;2�k�ݲ�P+:@�vj��F�pp^�I���{l����H\��Ɉ�Q��ވ#�\����E�b_#HU�u��"���z�8�a~�b:�c��容�	15�J�Y��dc_E��l���o\nD	4�'e�67{��7X��P)GfoR��P����W�ʾ�g�*+�H����C��xP�7R����l[C\ɷ�!"�У��c3@�tH���O��&��Џ[,JG���T�P���Я.h�F,}|���>ɏWM��iG~��A^�<�Ё~́TgU���t�@��${�(�t��:c�q�~��.�����j�������*�����&�Ü�cF0e�D˹Pm����������Ai��{�;�ցrT9u-�~��%�k��r�s�P�4�m�z��XHkZ-
��\ T�fvG�H>��� ��.�n���E��1�D�]ZU�&&Z<��Z[��Iw���G���L,���}{��=��=|���FF��w��6(�R*U����O���9�K��s�A�+
\�A��e��ʹB]߭?����������1:���>$U 5��5�ys�uU����z��E���V�"jc�Q����:m[�����:�v���G�<[�tW��K�&�(���R�Y0�bӝ���n��c��a�[��j@m�L�];�l�~�af  ����Uc1x���!n��k�6	�6!`a�����ZrӶC��V��� ���5����B����n�R�RI=�s��d��i�&d��q��?����Oaz��d�t�>b�]�v���.Ϡ���\�Y�w��'iꆝ+8O2���H]�(;r�z���;�!�ɵ�ζ�>���r��iP7�qؖP�`cVy���Sq���Q�2���~�B�
,^^�2�Q�b��h�C�ks|�ķ���W�Go�J��1�&���-�ѝQp�����v��������ߓ��>���PzV��������f���V��{��.�B�dZq�֦l���7���b�r�{3�LLO��KĈ�4L5Du��a� ��<�oA�l3�����5�5�X�
,ԜVI�j�Q-�F����h���+|�n8_r&�Xc*�T�r.My;H���յ�q�B��S���u7�]{� ��g�]ܨ������Ty�XSYV�Ƥ֙~���"� �I��|�]�5�Jd|��\v�|��"+m�`�B�~��=����(ٜv�_���\p�Eoθ��"˨���6��q(���\�.���G9M��!�u���|2��\���;�1H�Z	8�̰�d�=�=]���T��:��3�[��#fO�7�95�V�I3�5���OT�H1�M ��=������q##��y�P��݀F3��K/���
%bn�ee�u�I�3��.O��'�K�om�5	;S��ȴ����g͌��͡�k�V�A���V<��Rܹ����&g%48��*)@__l��	x62166�HLj�vͲ��>@P߸E/uɋ�C�1/?d���31�G'���=��MMM%,5Z��G9�Ԛ�}w@��CK4U��]�jf|�l��H1t��)*��<�=�z~��^�a/��3���<s�ץn�.}�]���[�m��t`�눢}�|����q��_s�Y�������(�?�h�K�/ţyJ����wZ�� x#�vF�J
]�D��3'wAW�S�Q�ݝ�$%��㇡1�_�����ùJe*��&�Q�������[xC��X�54���\|�4��5�Hk��o�����`�"q�dҶ�z�v���M����s��Ʒ�@����H��\�cW�:��`�����n漘����̼1�F��9�J�F�APb���B��(\�۠�?�
�(Г�q�i��u[F!�|q�F��U!#惒{h�b�l���k+��k����n9�����+�_�{ZP4'׀� m	��^gggЗ��������]��D�5/f�I���8�����焾�A��g�򿵿ǆU��Qsݾ}��Y���F�0�Q����o)�7BPs��o~�r�º� ~�m��0nj܊r�/�ڥ�f^ݤġ��kΥ��]t�`TY1Dr�mG3�Z��?��}yL_^~�J�d	{�uRڪJ� (\���.D�8]��:!��(~�s�w��}<'���fJ�6�К���� `MLJ����\Y�j�Pz��6a_�0�hsI[MPo�U��"�k�G� ��h��m?�u���]��';v]"���!<H��阜���'hb��ͱ
��x8/�v_��=�����@@�����.�BP$kI��������u�R�Z=+'W��+�RC�D�q%�|�C�hd��� 
�*75j�3�h��xA���T$�n��7��иy�{WQ,�v�I��S��(�wt�H9��2ց ś6���*r��-��O�����W�dC��ԫc���B��/D��<��bz�z̬�;A���ce6�M��Q9����W�]�h/��g�#ƌ���hh�]��֫�I-q]jb)��J�T3��2/��>ƴ�Zg^'˩�]�Ð?j��Y������lH#7���(��<�3��#d"�88�H��t+wW��~�dd�sh���fd�#��|����b��AWH0�����ݴ9[x1��'蕎��N�+�:�.��:�������"�j����g/L��n;�NMF��Dyi5!e���Ԓ��Jlγ=�*R0�^񯥥�*˭�Kr5HS+F}՜-;�k9T�-Z�_�V����&xPH7_�1��8|�]���-���g��m���u���Yp2�����������c?�뻺�)��P$.���Ľڔ�h�?mQ>�>S����D_0�-����s5�<���+��(:�h��7�ۍ%�>������:���$ɒ%��X�De,e솲U��!��B�}��,c����{?�s�9�y���u��>wa`8=j��yGU��##�q'��{�?5+kx<��8�(�I�}��wy#���&�^	�qW���I��_�����2GSC��C��m}&mnf���	8����%-�.��.@���Q�����"�|�4���u���-3xu���8���WN" �03�,��d���~ ���\ ��7��|���?MÌSuq>�� v�\����|JЖ�eF�S�]^������e���ǐ9��lA��<pR�?�7��`���\Ŵ��J&���Z_�Ǭ�� ��c�G�lS��j�������Z��	�,��.�hFJw��&���)�Z��b�v��W���������<��V��
��7�i�RC]���f{�9��Z��85�O���mڶ�d� ��Uf&���n�󟝙�Vt��ы��sJ˾*$&6�"��7G{��C���ӑ'5���Іlj�@�F�����/_����>�>Z�=�y祍=|�}�7���Ŏ@�F�x}�t�.uN��ԙ:G�ѢJ��[�k;��qp�� %��+L5�8V�૧C���!�m�L'?�0�u�O]��{]�x�����W�F�7��rO�;?\|r���H��e��s�&PJX �lW�F��n���������{BZD��Yټ0��w��W�^����q��bE�=��a�;��57�:6
��	�oNzN�'�ox[Rof���V�Ü���g��cF�J,Å�掕hf�-t�h��8k2b���b�"i�����B��F)xx��I�@�ٔ�y��7�X���/\)ǵr�]�HV�ـ��2n�x��0^�sB}S��񤺖1�Wރ�����%�::M�9�ɩ��ŋ.{d�#@��C�5a������x�T��S�a��.�-}r��k�~x��e���� � s��{��crbs�v�tl�.�=����]��;Nc��'����US������ɓI�.{r������f�n9�X�{��Kk��Ŏ}1���#?}�L���f�.U�D}!���d��ra}��}4�p�����c�vH�g4��&� ���V�0��A�f��������d�~��ܺc�>�7��X|���^�|Ț��]ϚBVBb�rb_`�����-�4�V�ɑ���mm��}+M�{��U���5�>����*�]�
c���>r{��Y_��:I���ܪ��O�߼hj2I�XOj*�ڏz���t�TN%�Db'v#�x���e��y c$��+�C?v}�[�5߉Zͼ\����
:�B6�O6b:b�'���;��"S��ӀX�b�[/ab���'�y�4w|B����-M$,%�B�E��,.�2����:ِ:����v8��Y���5տ������+�[*���:��0� #7�����BȘ�7\��u�HF�s�n��zݮ؝;'U(Zy]�G @����s�eq�w����{=M��c��}4�9�(h�%��u/��Z;�[jtcFGGǄ4����ڤ	���1��N9������鲇��'&oryՈ��� �+)L���,��mu�r&Z��b�M�p&xá��)~���}����/�P@qem���2Qy��%�D�ӭ7�8�������i�+K�� �˟#O����}�3_K񶵠�K�B�
�n4�u��m�c�_��9�OS	mQ�¢�����G��nn��k�{=�-*�F��Dc6��s�[BR�e�p-�C��J��MU�)��X�;Q��(����uK�eWne�ȷg�۷�<�
�~!=�V��ֆ+, BE����2��D�>��{�{�-��q���oX�ٰiw�������j_�%�d,>���B�\<Q&��vԶ��˥%��i�v5��j�۝����!Z�z�L�o��V�"S��Ħ?�����l�w��-�nk� ����x��߾�&�$��Uߡ�E�����{�l\̽��
/'��| L��O��*+�f�Xr"?��J6�4��.���,�&{$s6�nl̢�/NѰ_�J�ۗ$����֤��,l���~��z6�|r�((]#l��<�,��m}
 ����N�Lg��n�S�\]�z;�T|k�F���n;���<���6�=�Ss�������S'��~�X��)�Z��)ҪN��|S�]%���u��k=��|uTҞ,�=��D���VmGң�3��9m���/ހ.��쩖n->���mn��>��r���.�'�0�C���~;:�h^feC$����T�:l��8�s�J�W
�]]�;�[�'���P]3�f�i�֭������VA���@�ҖSbYt�m�t�����~���.��G���r���-���1�%�9C���>kH�A{cTQ�)h�)��mmw�*�:����&�����e�d>r	-bY�0
��{��S?`�?KTat^rY�ItG�/�>8�e��LS���g<+*|'�iT�+ڝd���8��)��n���戂rlS,[�'���̑ ;�BZ��E����ͽÅ܍�a��y��Сy��3n9�?=cRC9ފ��v4�p��(��(���#�r ����t1{��w��-���ʋ��@��4MD�j�@���]uq�=�5z��k0�2�~{�rEׄ�k��z��%�S�#�i�Rc�����ѿ����$��+���w!��&��>��Ա��+rGs�Z3�����vٛ�H�$%-!"PuJE��V���6@���j��s��U��iN���l�)C�ߖ�ț��O^	[}�����7����Q�nk�)���e���מ����sq��[v�Hn�+�N�%��z���Wh�ٶ�����^P��C�.-�*j(=WX`�16��2x.�@*�y�bKmbz�Y�Ct�}dTTk�W;�H�s�5���	*���?��<|�<8w�rJIWŇ����� ��-��
<��S�S$c;�����}� �6����<~�x���K�����s}�&��ԃ��]��bT�7Y@�|Klh���?`��]<��I�'�a���j����5�Y��q�P�1������H�Gu��zm��V�E�o��U���<����~����}�Kw�n�e��F[�ʫ�2�b 	�4�
y��j�0sKh��(k(x��p�{��!o��z)῾�טű�Y�SN!/�}����|!9^L�y��F���%���Ř�6P�=,2m3E� �W<}�����dy����x�C��n�mkQ�x�u���&�\`KMC����k��F�_�I�r'&�界��/�ҕ%��5!�p@�s�9�y����)���zy�Y�ۏ��C=���rR��1�ٙ^K������i\'���b�H��dnpe��K����؊� �ܗʹI�d���3����ż�ܬg�W��0�s���/��n�v�O�&������e����V���gQ�y���5�m4���%�FF����w�_�X���|ҺOZ!Z�m��!D5f^
{g��dSy_�SH+%�dj����ﮭmU���+X�i�>���ARJ+�}�+}0�7M:��*0>��&���M��0�H��k�qg2{@��L�e�Y\��g���.բ�SR#������{/��;6''#i�*���I���\�p�6�dK��_/}�e|m?����A�9��ɱ5, �5�72l����25B� �L����o�͑%2j4V'V������=�j���������"%`O�Sa���_SS���	?�L�Ʌ>�R���۫�)����U�0y6��x�O�q��c��{��I�.��I�$,�{\2�w��gs����b����S��B����bf��*?J�40����W���q��ʳ�s9����߽X��6M/�58+-��6w��?�z:\OWw�� ��U	�`0����6xP���׊}��0v�is��$iH>8�𝭾L�<�_�iSS���a����|�X0�����3?6u�R�8(��Gp����;
Pr�ӿ�XY>����H�h� �Ъ���N�������Uo�a��,�ׯ_8P�����7��]�y|���������K����u���9Y=9�����)�~�D!�����Q�W�u�v\臧w����`#�k��U�U��
��!�m�'}��[�}���㝦�r��w^g�}�Lư��/��)�8O�~�3ڏ/k�4_���W7L�Ml�U��OE�K�W<���$�Pt{w�?vw���5��Ս���?2�T�����|졅sk��c}�pM��+�w�mN.o��=�E��㥌t��iu��<<UP�z��o�0 ����{u������qAA��Oq%\`��"��_��+,_Z��4���Oa�80p����v7�����Y"b�1;�'G;-?�?UPP�"Pv���KR����'/CZ�ܭ׳��y��yS���_�y���Vv! Kә?�������\݋ze
U�yM?�ĳй������Y^�6OE�C�~I�,Iut��xZ֤[�l `�l�����'�q}�F_����C�Hj�v�	�I���l�58I�0�aLHL1��fax͖a��tL����Jm]��� 8k��6g�d��Nf��]v�-��C�[��T�1=�
��p�w�x�	����-c����"[|'v���n�HŬ��y�٤��6�L��.*Q�O�L��}Yއpqt<�8�*��/�'�g�ke�'}_!bbo�D��3ltt�]f�p"�|2z��O:^Gж�;��Y� �W����Ms?	;�E�=���d�EqQ���[Q�4���EDz�a(S��f�e�X-�i��r�� ��~������vT�|�y��f�{�'�]m%P����٢3>ME���Y��n�j7�[{�v}�aao��z�������v����Z�w������S{ǌ�;��r/�[�=~M��{��V䦼s�� ��.��
`ן�A��:=��-�S
�|CyB��V_�����Vx�%Z�DJ��/���R$�?<�?�h��e�UZF��x_�HZӄ��V�/u3[���R�K_4��Q~o��f��P�1���xñ��5i%?��mد�����*kW�]!-��^.�9��3D��I=s�zt�n��}ɣ�?���>����I��#�)���xU�r϶Aڊ��6J�;[A��l�釁������V9z/I8���cs�	�Gc�Ά���,�C���������­O��5K^��uV������1�T&[$�>t@��ebR$#�c�^ptpd�v�Ǐ�U��Z�j����I�ݺ��L�Ķ(X}-�cg���di�0�0갯��c����M���U)������g�ח�IPn���wwv�o蚡VK 6v����Ӡ�����GjKȇTA|^FP�UJ�]'B�h*�Kx��Qm�1@�!�ށj��pqC( !oI�L�)�=���Kʷ�NvER�@H_�"M5�J� R#섫FҤe�_���D y4w�����#L� wgk+�~]w�a$�#�J%��L+�}�܏�ӵJ�0E3�!��zrAbIJ��N���K�=�^�;�w���	�8R�}#�>[��7��t�c�� J�|�)&p���� 8A���k�`���Ԕ��5�ç���"X������5��*�Uv!驣��A�򾛤��[H˸@B��i���"��Rc�ϵ8ʎ�v��������t�{�����90�ǫ�w��`T�Jӛa�K���/�5�|��Z��8���q�K �ת�����o�U�/{��F��<8����y�����:C���������վg�m�2�VG%NًZj�63����~O�:�V�^�%�6p@C<�	�:����3(����KxvPm4,)#+�ݛa�`#E���
'�ֆ���"�V��G�ʒ#=N�$�����A����&��|��sլE��l:�?���Ffl�\�p��������I�	B$�;˽n/���֍3�HxGyw���!��C�]\hH`���<����z�z��0�ץ�$+V	�^���{@"G���d�ށg$�̈́>��鞓S�0:��*�Ìx>����dD�� kU1�H�$^�P�c�\K�yYGQn�hC��]��1lں" �A~
�}.�T�e�+�a�!����Tp���|f�)�Uqn}�
��\A �;�:���Ã�����ڴ��TW�3��-qe�n��%9\41�*z�@��;/�]F��u ﵽ�q����S������^`| ߔ!�� ������"�1��g��B�� ��SR�M;S�5���U|W2*���&�;E�$ y�Q8 ]�� ��%�}�aq��7<�"�"~Y��Щ��C��}'AXK�z��IL�N��:]	8���
��w	&`�����aF5ćR)�H]o"QZY�F�Dz�KF�3PjV�l:�	tq 9�7�j���50ď~D������p�\6�"/��弥XM8��I�s���ZT*�q� ��4��,�{橹����rx�^R� ��m)b�e�_h�vO����fֶ����(���P�_͕�潸2Br�d�U�3�.�����*���.��]g����"� �#�|�q���o��*�=`�P��g`�q:�#���ŷ�Ġ�ZJtr �W�e2���K��� ��@�&zoi)Yp���RN�bݪ6)Mgi���]$�����Y��Y�����%�JH�J�`����t%DHE������mO$�
ͅw��ɳM�3�⍭l<��9ӵ麒��o2��z��^fU~��(A��ݻ����C�=�d�_'�rD%a�
q�]�3�f-Ap,g���S>$uƚ�J
�F���ʀ/�������渧 !G3΋Wh<�����Q��*��-�gXe1���Zu�0��W�#�Anh���l���OQ�� oo����:G�Ф���/,���+^sxY=]J�����ڂAv���Zs�:��~F��m��n�	o���Lu�Ӧ����ʯK|V�p����\rU
I)	���hH�K<�`�p%H��������7��Ӟ+��-����)�,"b�l�+9	�P��,W�q[V��*٘"!��Q?����9�I��_��H(��	�gOM2Bn�˕�c����EKzj�;lHZ������5\\H>��O����S�N|R*�&��r�#$ж�4�.� g��*�G0��p����6��C��$݈VT�?
��� #��c�J����d�$�)FP0��S@9B	*%Ze��!G�7g��NM-��邂����wk�^HZYWV��|/O5ޘ�Z�ۤ�ש*�6���o���z�@ۼ���ߘO����� �.A��!�w�?=6�0�KW�o��%#>,��'�ao��������
�.�4��ey1��s���B���M(��=�~�Cӽ �S:�7��℺����W"6�p��������1z_����~��g���]�I��R��zql�Ƥ��=wx�We�Ѧ�J%:�ŚB�c��C���?>�s�nm����zB@ʽK�=y�0��2d�p�S|�����������	�ل�p3��3P;:��9"(`
�B� 摩��Z� ���Ç���1;�ǫ}�Ϩ�C6�.��GC���$���D��i2�X��b�5�X@ ���}����lѝ/ʫ崒�J�R~溒���'OO]k��18e{	�~��D���È4 �a�AJ�G�w:��e8�L�*5ɕ�p*�(�ܽ��B�)�����n�BŒXχy�,]�Z,�hqF��B�f ��ކ���*H��; ��iz=fК_�GK�#	Xge����	��?��h<8j�� ���o�N��,��n��w�u�r���	����l�a�_��s-�� %�i���[��K%D��5��9��G}@E09K?�a��p?�d����x�'Dg!�b�w~�|�o��~�-��3��/|a�C�ٚ�I?�h���7��*��fe��U� ����{�Ԕ���`0��]=�*�:+�|����mn����'� �τ�G���m�ixwZX>1h��5�`���p�=��)9�h��g'Z+�D�V�� -�cb�r�Y�.-�� jn�)�t���9*����ԏ%���K��Y����Ea��ؙG��o��1fW�h��{�滿V,��KP��F����6.{v��`���T!��F'6k���ҁʏK&�4���o\7�]�C~�:��~��kuLJ�g{�n�膞�&d����[E Y4T��2Š��K��������h`QՓmU�Ԙ$ō��r���r��%9t͈�T���+E���rbU�0��y΀�֕��1O�s�	���مA��#�i��U�!-mN�Dí�k�[����߿x�^��@wCϚ 
gh` ъ���)o;�d�E��WBT��~��C�T�bC,1P�.sMnT�ݨ�?8�:��w�ob���R�n�NR��G����tЈ9�F1c�7<�ֈ-�ѻ����j�Sj�Qx���'ۉf/N���<cDJ��y<uuː�sL Պ�wrF�U0�G:�q5�q��<'�&��uR�#x\����ɝ^��2<�m�§)�J�ޫ�W��خ��u*l�2�T-�?3߫-`������6F}����x�Y��H����f�h����| 2x N��!+�4O%܇7�f�âQQQ��˷�g}���F���B��B�mI��.�+U�����x�M�4��_R�wGƯ͉7����@�<�-�����GjnOz@o�oŴF+�� ��t�;j�L͘��Y��N9u�+�|����b^�lm<l�/?j5�vGkjjV-
���q�,F5���lm�t$S�$�v���V��J���h0��_��ზ��9���+����9����Z_����_�s[~�aim3�io�^/LEFЖ�0����Hi�aw�ՓvN/ڔr��Y@2�[�D��L����`�Z�p��ެ.�?w0���Ƙ:��5��爩�ԽԼ�5G�8��x�4���e��һ�C���c*�����M[.���A�-0e׵�����3��!U4�xQ�������X�Տ��9r\���U�����ä*`����E�/pDX�)@YmЋ�Z��פH�V�U����W/�s�
;M_=ˌ�^a�F?����r�G���{�(((}��1�����=y�I3�ʇ����Ѳ�����Z�}r
K:sU���У�nh����A����+�Yy/A���u9����Y3�YQ�9J|��/����� s }��u�Ө6;Μ�WO����Fݩ�n�����Jf��%��	O[Z@�Zf��-.:Y&ǈ?˅��Ԩ	��	]?8���9���W���Ȯ�G�Ⱥ��7Gs�14c��v�t�vw�[QO�`���i,1�kp���L԰�64����-��]��BL�o���������v�iiO��.�֢S�w��iC�"�I@�S-�4t��u5u�(����)�i��քX�]b#��{�\����!��e�+�����(�#hS����"o�]'[�U?��keo+w�?��O���دH{}pz��!������^UU��Ir�Y�8
v.+[ z确���*@���)RgW��fZ�CU�+���'b����;;��o[<��4]雐�:D�)?S�j+��O�Q�Y��	�/Ǵ��x��s�{��[<1(��_�C~è���У���9e&!�$
�ʽ{���2n��֖ӵBd�������5�a�gV�T��l��^ۄ���£s�U�<>=H��O4�0q�$��]�36Q�[�:���Z�L=LE��� kt[���,A�h\�(6�w�%��_��C.|t(?�Pk�-x(H)VV`�oC1��8]�.cy��'<b����JW��� �5pXF')�ome�.��I�N��M{ۿ��Ol�e�b���M�N��Cx�k�DF��Q�]��iu:<N"��8Q���h@qu%'��0Z ��<�3v{�1f{en�X���+f�h������b�a���^@ ���I�9�����&~e�ܦj�����efjW��'�S���p�|���ɽ��d�����b��_&_~�Eu��yp@Z�o�~Y��! ��V_���1A��ψ�@�y��D� }�ׂWb[k�樆qe��d�����+����J{>�5���:y�r����&h���h�_�ō�Z�aø��t=����,k+�e*8PE��j����Q�[jEa�q����m�?]�ӌ���u�V�¶ҋ!M���TZ��0��4}2P��0J��R�BbR��Y`B�[,�=��m����ukx���7��O� �	�e_n���kfL�}M��������)j�-�X��t�^	�]��>����D�|Ft��j��.i9;9GLL�h���0!c����]Gp����3�8��S��՟�c����$���ݨ��q'Id'�������\��c)�`8T���]bkh�?_}F�`��y2�V���)`yi�����팓>}���@�z��J���8G�R�auc+Gg��̰��y���ԏ{Q1��8v���B�~����Y;e����K�P~���ɐk����h�!���l�TV���I �9�U!fy���XY�� ����i&�%��<�SX�]ҚM�C�n��ՏA������NG�O!��"�ϑg��P�9^���,&�<L�ﺉ	����K]�6�i#`�hs�!�����8x�Ѐr%r����1/���ޗ��2:���|�������@��$3
3���#梃����jR,s���ʥ����>?]<��Ly�/���*e���Asʀ����#(�ߏ�3��
xW�no� �M�A� 9��Uz�w9FT�[��+��|�YX�Q��8�V^e��x<��@��WD�q��H�p1���,���Y�$���p�ڻ��J ��O�9#Df����'�� �T;<3�2*����)�JrY�P���r1]����>�^'X"M��j�;�1�X	� 7]�D�G�g�9z}'�LO��^�&W������:K��f�f��C/�|�<^.͈�����Չܘ���P&�2V�-,|6����%�2F��y[�k�'��X��E[��͡��d�~�Rb�	���靰�)&��Ku��mkIJ��	:E��z��J�gG��)�	߄�,��0a\��:F-�_�<c��*�W�Gx��r�k	��`(�bG ��|]�9 W�=҅��;#�+�e���@xuV�9�z}���뿚�O!�ߢ��S���k�Ӣ���`Һ�\Mq3P���Z<j��Ў]���Z��#9?��<b�����4���RŌ�M�[F=�qv�i����1h+ʾ��� r;M��qFe���7����B�E�DC�H��Ø����=3�CىϚRV�bE[��2l�_4-����#�M�=��4����'+.U�Rz��'�M��r�#���O���役N��2�wgw��C�lD�2�-_���nx������?^q=.�O��� &�՘�1T�'TZ(��p�y�@>�6�=r���->�gu����%+U��\W�ܧ�p���|��o7��(�~ͭh�[9�j��h^R���6���x, ���i��ٓ�&,v_�!Ch.�ĩeXWr?�*� (� ^��=�+HҭG�&�BY�>#����,��TZ�:9�4��@K 1��u<gqͫ��2���%8+�s�T�?W���%T��Iu���5��-7�C��{�Á�|�!#�;;#9��O:���"�4����z�����������98:.���ٌ�)�a�L���;8�^��=Z�?_0���s������7Q�b�`��Ŏo�6UJ����}�����h�e
���CEEk'���lڷ#w�X5���s�.�@��|y����=�$�ʾ��%6�3�$h�v�B�����B�x'$�@�QM��N�ѐ>�T������Y!�%�r(*A7i_3��{�ۿs@��zs������� (���o�E�R o%�t~������ ,
򱞟Ü��fC���%���T��l`�B+9wR�_WY[,`�E�*a9�@���%������Nc���W�f��q�?\r���j�A? e`OE����|��&���\���5P�H��1����SN�n���s�����~֦3���ʴy�����9϶ �ۜ�(eL1e�\��~N3	\n�(#�_fh�V��&�J���Ď�I�ɷ[Z��h��iK�?��:Θ�=9b��Co�seaJf�P��0va����yIV���t��\JҌ5)��96��?{��"�9��jy��Ƴo��>��?�a�N�졭��o�_�ǂm���o��S9���F���B>&�p��p:��o�[b9����>45� ��i�һ�B"���z�]䇫�I�h��CtH¿��3�/���M��L����f8 5����~���5N���+��y�xP�ϒ�g��"��������
��8�ʃ|�P��vlۯ�s����C"��N�X��KJS�ՋH�d���)���s��z>AJ	�뒫Z���Q�J�iА�Iw�i�P�������qu�1:Y�Y�A�^j)�h�P�I����Q?����=ڡH<Ћ�Jݜ[X;\^���^[��Q�w�_ş`AR���'gr_)�8��Z��w�������&m�7��&3y������*Y�w.����n%n�F�݉��Ȯ�J%_���j����߭��z���M�c=��A��?!����/����[�׮^9�ZYگЏ>�ۤYD5O���썏�{U��fU_�z���bq�M
���K������4�'���r����7�P�&m��z�f[�lnz����~;�g���	���:P^��8��������B�u����H��_������_����F�a�3Q�e�RiH7<x����$�����W�m}�k���/˽F�li�G�@)Z�aQQW�e�W�����n>��S�2ˤ�\\&9V��oV���{XOdt[��c�^��8�٥5̪�p�:{~u 5ƩV���Ge�V��ۡ���ne:32���%b[�'��k��|KP84#���_�#��L��ٸ�h���=H ��c�k��8��p{/�\��Ү���Q�ᘎ3�OqQsbpc��X��eB_��������_㟆|����~��ߘKv��!4�0Cԏ�h��2 ��Ʌ�l7c>$�h��$E�3ͯ�յC�Ws�쯮?�������[>�C5!f�@dR0!�����r���6L?��F1��'�)��{IF�R�j��;1g
<
�4fS�Hs$j�`�|�a1Nmh����n�px.�F�%��f�s�I�ɐ2KRX�	����������֖�i�Z��6�T�|����jwҿ}�w��5�|^϶�rZ�%�ߕ��6ӾN�C�����a��IL<J3E��B�q˛3��m�1m�o���{�̩��`�2;�lU��?�ݾ�����Ӿ�U���L�g�������"h(h3�@��߄����X��q��1u�߱/�1a�	_���/���y��5�j�m���	qȖ
#`<=i���SS��m�r�:�y�[ۂW���6�K��V+mO�Y3�H�f�~��π��WB�r�_m�F<�Ty�y��� =��j�qK&4�v>7���9�� j}��Jr�'�fy������8L��5��Hr��PWAT�������p�iS�O��\J�ۘ���+������-U�}��;h�J���?SQ>����@� hV�}/���Bws��|&�"�%i�_�l&#�������0����hc�D��k��DVL�8k��o�T���O��o�l��8�\"Mt�)��0;A:����z`������1��I�4�T��XvO�V�sk� ��IK�V�NE�^���[!#���ѮT2�������d��ʪ0�^��I^W��!��u�N�q� 6f�����e�T ���<�*-��s����k ��AU��Aq.�l"]m_�+�kq�/S蹚tW��G|�E@;򦾫c�`�	�_��V�(�k�mkw��S��Ӳ���F�BD��Uu{g��e���y"K	{�D<��T����m��N�8ê�%YZ��o��6��F�l(�0�h#t�B��������c ��y��8�ԯ_�m0��]AظN#@x�]�.B�w�n�;C�N�O}�Ģs)Z`�b�AG��&MS�9����y��N<��ڪ���l�� �QӢ7Ѝ8;�����/+FDT.�j7��jWAX��Ł��Q���'�`�����I?ss��W�:)�J8 �g�P�͔X,�?U<��r!�fg{pt>
J�jN4�֪x�����k���Dje��~������7�O9�ۖ�r.
2�>Hۜ�����4�#h��҄
�Dc��,�Ӯ��05����B?
�������+�%o�)��m�J��a���<���ʷ�p�B���������	�cM�z�d�����c���#��a�����.W<�ǿ���R��/(�-Rxhsg�$<r=#ֺ�}<N��Q����;4H�։k=�u�Z�ƈ�y���6f�Vo�_ ���j��8�=�y�!�4.W��T(S���W��|\�P�����UyZab��\ �<u�O������iR�[U]��
��.�.�τO��te!�(¤~Db���+��yw�<�ݟ��#�[��f4L���7���d������IDt���)�Z�,,8
��E|��� ��[��ƀ[3m�˘����$H��Y[���&��B_��@�`�M=Q�> ����!�<��9�5���J� ��P3���Yu�*�Ma�����%���.�aD��eiP8�(�U%q��Z	'�h�b ���Ġ�SS߱��voE�p!�H�y��RFz�^tݸ"g������;'ۅ�Z���?�.b���h]P�r�ٿb=��`
D�蹩XN�)�t7q�a�"�׹����{�Έh ��.�P�Aw�x������  �Fǣ��ǘs�X.܆2�b��\��T�Ľɖ����9$G���\d�x�dr;AkZ�XtW7��>s�.J��"�
:�˥���;����k����������D#��L899]u�c|]`b�c21�jj^���*.)�aY+�{���;��׽r�;rgɴ����g���	�����r5���[�T�R[��2������4�}�b`�4V'X�m<د)���%��/��t��0TF/��\�w{1�upI7����(_��X�T���ܬwAfa��FZ�RPL
�^���k:5�Q�ښ[����V3����s�&?�?��	W�rƦ��J��na�J���<p&w�m�':6'��C��Fs|���?6���u�X�e%)�g^^w�4S�e�DNEҢ���������;qߔ�p<��,;�9�Yt~�Խ���f,sZ=n��m��Qm����!���'��� ~Wo(����/ɩ�|+vC��2D�?o����Y������̪����-C[�^�q}Kn�����Y۩/7�+"�-4�.u�8-�����b8�7�ʒ�+)Vu�T�؄�E`x��tY�׊�8�\��{͵^��R z8���ءa���yg�z*���X7�kmj��
��D6������'�˂���B�� Hغ0�2=#]\�D"b��v��>|�=�>�6�"? [Ď��6�)-=F��?,�m�HA�"bbb*�����|��	j%Z��J����n�e���j鋭���G�'��؛Q?�vY��S��6�fj|�~-���X\���B7�u)
�7{V��}1rKq�#���
]�I�s}j����C�i�ɧ���Z����"�^Ʌ�G~�ѨM��^\u��_t��<�sP�x��̜����T�ƹ�f����$?����%E�L�XDtL�T:~s��Epȸvy~.��Ǟ�׻a]��[���A�<�Sb)�>Mȝ~���b(�����r` Op�	D�a����ܶ��������8�s��2-a��!,Bs����4��e!���b�s)s�F�%��ۄL�{�i�2�~~���9����z=�y|^㉕�QU����	uuu@ѤGi=w���<�Iv6�����TttJ���?��G�0P� ��bK]�[Y�,�c�?��oee���g����C&��-��������F�>�w7��'r��w���w��g:7Y�Q�&��yhߣQ�X����I}���v�VU�� �c!4l���S;��ɽ��^@��c�MG�7#9DS*���0\$Ŷv�t���� �T�d�_El�'u�oo���WP�<Qp<�­�yͼp<� �(����#p �e�w���a��/�.t'�썤�$zj�o��yN%�`&�Rwc�tLB�®�	
��ت^�&���;�f˜��sG�:�L˹o�Ӈ�j>�N?���l�����f�vR1���D2C&�Fg̀b�״�g�	���$~�+�l�}n|�^#�3�	�Oe/2'���a�aF���UF�w���=-�����p�4��)G-U`�`�a�/N�;��J�ރT�fǳ�qoOYM�O���>b~���[�8a	qY�(j�Q�-�W��M
OQMLL\���J���}t�����>��.��zf+\g��ya�N�c��
���K�kG�qUk@Jp@�<�m5� ����,�=�1�~���,W$$�Nh�ێ���À=��AGM7�ABlA�A�ޟ����oa���1�&)~=�Y!��\j���sx�w��[z��8%�����p��ummm��n�Ñ�ߵ���=�c�=���h8�e{� �>O,�3B�U��J����Y������vΏ���c������=y|*��H�MɁG3J	g�R观��|~� ��N��h�N�ê~�0��)�4&�Mc�ǆ��L�gmV�	Q����4x.Y��5;��l�ԝCTZ��=��>	V%p�{l.�!�_C�������x`Q�[�lQ�M>g\��	Q �r��o��s�<���[p�6+�0�(�����KS��o���俭�ܯGn.�2���<F��]���ct9�A�+���}��	����~f�&�\��^��zo��L�	N��>����P�%!��7����_�����A��,�zO�x�_ڨ��'$�@����{Ԑ�s�5ů$gw����$U���s��}�?�,�L ��=�5E�8�ͱ&�-�(�<7}�5!G�hU�W���{���s��M�^cN�|RM	��?w+�gk^���bù�D�e������s˫Zq"��<䱑G>1D�C8O����4T�C Rq:���O����B۬�ȇs3���>��{��Y��!*p7�{&Y	0ߣJxkE�t�o¹�����f� 쨪��g Ƃ�����;(��-���2W?tН�#�/NL�⤛{���s���h�.>�8ҸڪP�N��a��NFNIa	pgRJ�)n��?묭U�Υ�D�	\��M:�=pɑ �C��k���^��IR-������}!>���I��uΞ�I*/���ۿ�K��/ɔ|�����n�B'�&G�^?�%Q��#�CA|A�iY~b�QRU��4r���8y��s�D���[�G�
^���S]�h .P�@����[�T����*S!n�(Y��_9�75�~��Z���X���S�k=#�ױ�7o��/a��#2�\k[i1��ʾTJ�Q櫙]��"���83z���s��3��)a nB:�Q��hǡ���_�e�bo`�U�m�ȷ��!���<�pC�;a k��Fq�`�%�P��1�w��9���5d�>5S�P-3����ĭ�JE���(��3Qr�H@F�Kx"B@jj�q� � iNg�_���l��LPa�/��B&�)Sׄ�������R�o����c��so�#J�X&�k�AK8a$r�֐��E����i�I\283ca㟸��X��*1N|�Q��S�b�o���>�K�y�P�L)i�Ik�h��ũ8�d�A����ݟ�X��t�� ��s��+P,�e3X#�T�t�KMM}PDe��LV�@MQ0C876 ���q~��Ӣ�}����i�?�h�ͺ.��a"�Y�� �7��K��B�r������lM����X;��m�aIx`���OL&<N����B�.Y�I88���箇We����9YB�O@������3�4��4����ct.� ��Q��Ca��]%c|9�Ǣi�/�>}ز9�4��/��U5uˣ�?��eE^V�M6���v���`<��׌l(ݝ��}/�8��I3���z��&��ȃ�/S����j2�R��Sޏ� rz�5�j����y��5���n�Wc���H���IY�N��u3���$�a�B<�M(���Y���\��C���f^C`T�
,6J�#��v_�|KL��j��]
WkD��v$��FAP���Yø|L����U�%'	=$��+��1��J����j�,<��n-����qW�y���f9����;��Ǹ�ʪ2$�/���z�!?���@�����߶_�Xv'������Ț�oU������V"����^�%}�S�m#S�w1����c��TSm���z-q��c�>LyD*-SܜB�7v�R*�L��"��x6ZUQ���ڊ�L�C� �G�ܛԴ��+lk��9�9�����oQ������8�4�س7�|�F���V5�Yl�rܓ��}1�CD�ޙĂ9N�W�����$Ci�"V��X~~�˸v����J�wc�90(̣^|_
k��<�:i���P[w�䠔�K��$U��|��{z�����X�����U"OQ���u6����� �Z!��B}� �j Dss���!;�x���6.��猻��<��R;�M��De.xT��˜u�� G�_�uB�����q����yA���9�Q��#~�S��V��~zq�zcg��3��x ���xie�QW�y�l[?����H
�0�Lp ���%{G,��J<>g^�'l������E��N����/�I���ޮ�'�A�o�M*���̖�Պa��3#�;�������u���ujc}���|��4�81��i1V�^���p�x�������j�U��iM���W��#׆�HZ��x���݃�Q���Ta_Z��)�y��B��@��3�s��θ]�G���OC��{sZY�eN�C`��k��ٌ`��c�H����BӺC�7��۴8�@�������aOk�|��>��O���(�T�l�Q��� ���=�.s�O��_! ;1����/�	�B��8��qB���D}wTgY�={{��e9f�����|���0��D8>����ΤPAn���cN�J�������W��z�-vo:WS��n�}�x�/���M�L�޳��$�m}�HvQ���s6�$�ծ8�G��j2R��:%N��u���"�fy�� a�R �KT	$�o��4�
��}�a���9�"�� ���� �tA.GE�Ɂ�{�c��Jѡ�7�N<W��q��_#j�O�{��;r��J��O�͛7�5�MM�����?�p���QI�Zߵ5�:isKo��X����3A�Ӻ ����������k=�Ʈ$)�MHw������T��;%��=X����՗D���c3e�� �:�ˬ�?�tz�w-7���~Ommm=��������h���ZH��'���;3�Q���8���ma~8^���	�����d�kv"�l�i����֩g�=�:X`�v�ɔ?���Ҙ"ݙB��o.��lU��i*{Tˎ����3��AJ�R��n��*���,Ѡ~R0#��|0�W��o���SX��j��c���V&D�Z�^yU�3�3�%�Ɵ��,c���o��`J~��{36d�J���&//!	 ϋ�vbIg�Q�r�@�nejgm,X��K���I8`{����x\`T��7�M>����|���,s���=�����-��6���y���R��'��54r����<I���'������9@�>���A%����a�O���/i�c�8���
>JSw�&p��g#�p�F�r!�	x�3�QU��"�pa:��'BKU	�R�*L��.�N?�U���˺����e"7`�����b�檱�D �x>V�gw�A�"��Zu���롦Ax7�D����=7�i�to�Ox�N7���*�.}�)m;;��B[Zq�U?@~�����>o�waͯ�<o�79w�Fl��ޛ\�;c�q
�<������a��y|��v�
U^���������`������hH�|�+�=����/F���e���<��H J�	�M�9J��m'o���5���&[�c���o�����U�Ё����_>e0�����T����H.3ʙ�Z1�-�s��{��z���5w��	p�/����3�7RGŕ�V�X?s)��t/�J�h�sK�]2P���VO8�ڂ~=�!�Z��}ȹ�D�2���k�������;l�͒}��w���JX^�k�-��T@����6��)�Vu�p�Bg���yU���c �����˗??2�;�|�0���E����9$�ʡ���aVUS2��3�z>k�-ů��.S�F����N�Է��h9ReK�Bkg���c�px�O���JW�,n�k�L��cH����N|��ܻ/�N�˻���r4RCP<�ր�@�_��D~n�����nKG;�Gb�<�ƋB>0��Ia� ��e��u40�!�t�9�NkS>j؞б���m�O���Z��;�#}�-�2��.i]:�Ik��0 �74��e����o��z7N���Y)D�*0���_�����[�&#��pnC�)A=�U�ḇ���.,��k�^~ۇx���:��⻼2r̂)N���5�U'�d�ET��$��踱9����*���E8�D{��7m$�@�����Ęih�; �h���ǅ�17=#�-3�6��㡖��M:���8�	 ϫ����F�f�3���X�I�m%}��e#ԫ���;A-�p'�g`����S��S)#`��KOL���u؝�>�[�81�+��"�,C�8�?���k0�'*�	k�i����r�r +M$�g"x(�õ��c�>@N�VM�����Fɡ�	�/I}9�¨��4�������u|]QO�@����c��� O;�V���sDDE��ܖ���T�J��FP{Z�����S��nm���Ͳ\k�K�,�/����*ON6z��>�bȩt�g���A^i��P�qQ=.�+�����`Ӊe�;��X�)1��'����ϝ��xY��/��� ��k������kt	����¦�Ao�8V��C����Q����l����*�C8!���(!�U7�1f�#! [��F�4�#'*O� 2z4V���D<�&��PXj���|IQ��nClq"��|��7�)�z���� jq#��ͭWc�,x�Q2���	���Q����(5x��V�>�]�о�a@�<i�'��g��}������p>�� �:���'����o؁�씟��L�
�(/0_�ژ��)��A�8��#�Vx;��f	"���-,�\3�~(,�&-]g��A`E
�6P���"�K�g�����&�4)*&fHUߋ���2�������/��&��TIpWu��9oa��g:ۈ���C�Yr���ʇN� �t"��%T�8~�j`��Պ�
�V<Qd�|���h����z�tA0Q�jC��M�O�K�<njJ�n�t�ԶҜ��,A+�;r�$��J�䯫�o9�o�<��.����% ��%~~�;dO4R �f �����+k͉�KccA-v�g4�v����^����_hM�m�Ń��&GvEu���R���I�73n����W�
�D�#5�� �������^�9��>�]�T<��Jk��)dA-�D����_�������Q �MkD!  �2���~h�B���F���8Ӭ��,3��Ь�3J`��_/�ݮ+�+�*��u^#�	p���G�y�2\����ʉ�C/��1�K"�BH�g�>T�����O��Q�p/�`�3��u�͜f��x`+]c��.�5P����	tP���m������
$��9r�</xB�1T��3�p�|��X��[1K y5�S \�) �h��w\rz�F��:�6ۿi��\"�ܒ�t�-��=��">z� �H��)j�Zݍ�����d��бDߚ��L'��_�v���08ul}}wwwrrrd�i�g�rn�m((É#9���!�"��橂�D��Sx������QUmI�������Z��a��F�
���W�ׄ3W���\������5n^.l<�܃e������m�i��;�k�U�L�����5�$J �k T���sQ���q-6v�����Ő���eeeo���Z*��'���Lj�I�E��̃�@]CZY��(����42��:	�7�x�_���$�F�����鍍�!]�u�A��(�O+�{P�Ӌ���2R���MO�/���M��9���4x1]�c��j��M
F�I6�����_;����)+�s��+'�9O4���S�X�AP6�$g���$��-4��:�|�6[@*�V��}�&Wǌ?�)����|'�"�%7i�Å����IH���K��v~�w<R��TG�#��<�f��ElK�#U�@\&�n�uP
��U"PFhe�okB_%�h�X'}�?�}�$�4S +i�U����6�g,^��H�le�.� ƋJ���r�\H�TUc����,x�(�.������/��{έ_3X�%h���s�,���6�# ���sa++��
H����������{�2s_7�5�����.��\�啧 �!r��de���Vd�z>��|�B�lé%4b�ߛS�Ğ������wb^]4��h�jz���9��w>���7�K{7�l#��:�C��PD^4C@κ!Ϭ��_�K~y~�4C���I�Z�̾bo *����-f�«���i����9܆�Q����
�#��
q�T8ۋ��ǁ�Cd�Kgގ����5��L�wۮ2Q��)opl��D;jk��h�f�����8W��{r��F��f�q"�U����vcv�*Ph�3�,R�ޓ#|���I�[�p�y�|q��7��8^ަ��Ad�u��.�w-�,P�4��舱@ܯO���R�h�(�f!�f�v҃Ĺ}�C�3hw,�Ĵ����~�-���[f����5~�������9���%ݫ�}J/��&�^mS�[���X���sxoѬ��1~P�j������r�l��Y�8�͛�~jw��7x��k�Z��'���JR��:�J��������Il���E��'��>��`�F?��ωW3ÃX�Z� �gR�MU������ܟ�]�����Hu9�	5���~���ƕz�=;�:8�?P�Қ���h�����Qb]�v�Muuu��~5Z�Q��������Ė(�USG-���1�Y��Z>%_9e�,p���&V�jz?+�u�}�! ���
k��$�;}�o�ņo� O�2pd*�y��f�!z���'���@gj���e6R��Q����:N794���ѥ����`ײ�3<��Ҷ�-}p䡶�k�c0�sihkX{omi0����Y�g�\wV�'��a���ʭ��[������6{\�㭜j��Jk�{�8�dx���j��I��Ne=��B7��f%�&�Ρ�m��Q<z��B��ɶ!�� ��\���k ]j��]T1�>����o2TL&�g{t&��q��}�u�����_�5�?條����=_g�	ku�g��HN|�������4��0�/6�{#��e��-�$���ެ(p�ͬJ]	Y��[+o�~X��޷�y�\k�u�d���5pd?��� �"pM7�'��ϟ�t&କ7iP9w�P�)���[�x~��� ��^bC�L���|�w�R�F�U ������	Et[
E=fx���~c,O7�-/��z�?3V!	H׸¾��<�j�Řj]5�y|�Z)���Ě���%�Nb��L�*3[sRˏ9�5h�=�	9/��9� $��|P5�w"@��c�$�7��ދ骏k��>$�F�x����c:���ظ�0��,����b"NF0vN�����Y��}#�)>��f�6�ET�H̾�ʅ+�?�=л�%�u��D�Z��H���tD�TEJ�$m.b��MR|	�[sL�9Ud���K�Hc�=gW����'�����.A��9YP��ɝ�N�\��7&��.IW��3�S��<���x��^)#����Pi.ޡ�7��W�}eq=}q(F��H��� 6�u̙&��oA�~��~T?͆�T	+�v��W=�Md���2�y�A�/�4{��4�nY}a,�f!�zR��ߍ���y
Ԝ����⎇�z��0czp�Z��s����OXD]S����w�Fi��W��b��UL�������$���w����8%š)w���SΊKR��'b���Ih~S9l+$	Ԧ�)*��/n��j@<O�#VLi��&@����@���r��x/�8�o����w3����~��ӳ$�w:	 ��\��;*<_���k}���aB�U&/O�l����E�^�|P;S����^Y��U����Ӝj�üX��u��S�2z��}���Y�S�?
q�4H.Gc� 9��}��ıU (��O^���>�Mn�OP�"ޓ���TGe*���_@Y�4��|�O0�뻖�����Q�y�8��-��D�2[��߿���n�?g9��QK�ؿ0��.yWl���ƹ*r�آ �e������,h�K
˱e�n �SPQ9�|ӻ����vx�O����K�֗�1�--h�l�o�c:������W -1��p�m�O\G=���9���WV�[(O�nK��V1��Wg�E�B��%���BvV�W|��+ET��@ۊ|����͕з��P~�L�\tG�T4��部w���UHT_�@�[��T�\g3Ah>�����Ϲ]��b�ϙ�ם��#���!F�\����f�������!�V��5�IIOܱ��7�,#�:�.6W�?��S^�~kA�L_�F��&Aɋ��>�uhl^G�~ɨ?�Md�W���n���Ax	`qf3_l����D,ǛH��3 �!�
�l$��XGl;��Ԅ>�FS��F�~k�3@�ԗ�4�&Sd��I�� 3�mm��Ȥ�;�_&P�>vS���g�K=�U��ш^�$���邸�ት�w�l�e R�L����}�+3�4�}ѐ�59�(k1uX$�e�FF�婤�_02{s���S�mZ�)��w�y$?3��PK�R��r���3q/�N�e�6ڙ�5�����է@�J,A���[�C�gs'�`���=_Q>0p���v�1��:��( �e��A���`�6��r���ޱ]�1<:驉���s�����Ň�b8$] ���i<	:e�
�7ܱ�9*ֱ.!T��W+��^M�M<�;�7�4fX�X۸w
I���К�N�+S���b�qMf:Ě��I�����P�)ʜo����CrJ?�A<��9�~1�=�@;������?���;�l-S^��/0�C�l�A�D2[�!�g�$�h��a�0h���nVCL���ˡ��bn9*t
ִ6x�Ñ0��V���hFHZ;�je�}�k�� �?�}�I��s�������3��9z�PP+J1�p��V"��i��,�=���/CC)B�-38���h�t]���(�!�Y)�]!F����g��#��V.���'�����l�)�E�W?��Ŭ�O��~�����c���D�Ļ���dQ�Ʃ�ӷ�!J��~�eH����nA�������۝F]�J~�K}6dc���WTF��߾ǈ����(�z�z�#Q�ߎ���޶K�N�_�b�d��I�Œ4�?��Pq/o���m�xu"jA��[����+	�/�iq��%�KZ���ucա�<h���v���>^y_oJFaU�B���sKk �+3�8��T�
��Ό��9�R�L�4̐�1�RR)cȿ����q��Ի)��U��>�~�>Xޣ(\��N|I/BS�1w���;ф�-��Qt���6:���������Y�}a�����M+���'��"�g�_Iа[9w�ܡ���U�.!�����e7x���'�@�j9U;5�A*����'hE=z�g���'�����n��'�n2q���(�B�k,�ڄ�;@'�U+x �<���ѽ�~W�����g"�٘�ΪV�~?��}hJ�U��
��I�<^r�ז�,��h�
�W'�jQ�?X��>���?5N��_�ԿxA�ԣ�r����1�3o�����ڟ������`��G#��}�h/]�S��n����.N��0H�(���J��S��-R�r@k;��RS��x�7�Z�B�	?`!}z��*��j'��w|iz���M���*����N�?�����ᬬ}V��	& SR��\D�
8�
S���!YzS�f��@� ��d��h4ö6
#��p�j���(>��GEF5�1y����3x&���Թ�+CU�k���y�F[%�*(��w]�O��t�&�/��y��R6��Out����8'n���x)��LHF!�4]��0���@3�����ןd�4?���ͱ�n[[ �=(E\��͔�q�߳1_���25@΋W�-�wobn���ѱ�~~G/��9Hi�r�Iǃ���~y�[H?�L�P��M�H��^�h��+�F�l�,~���__[���4���\�Y�H����v���p*h"xj��7��W���jo4Cٳ���!���߂���eOz���>��a2����~E��R3ң=�m��!y
�lƥ_�457sp��U%��~�"~H���o�f�q�����	��檏��[

Ka��T"��y�Q���M�E��	ϵCU�II_�&�lnyE��J�Ǜ%�v�o����Mڙ����$m��
#�����y ���H#����DWt��Qf(/��צ��.V:��<�����e���~��vzg�J�Ձ%b��p'����Aɰrf�W�5�5^������ϛ�o=�/GzNŞs��ո3y .���~�ay�C��T~����amTP	���V�nw����Z�y(�+t�@�ݗ8���{7��:��qY^Y�p_ɉ�)�E} ���+�	&T��|����h�x;��G�`����(���x���(Gq�<�=,���otȭץ�(č'�\����>F�9~�`~ݎ���6N���s��nhg�W"��4�@�W����	1�<�]��`L�I߂�"y�?ޞɓ����@��E��/��@�����I��R�<����J=�w����lmXj�@�6���U�G��Z�>X��
RN�#�/q"�敲s�h��Ù2�oZ����B�e(^$L�G�:l�8i\�+}�.PW����tht�@$t�dt��}�9굦�� X;|[��(B��9�x�(�0����B�{eyP�(��� ��L�E_�+��ks3��1(ڋ3 +��>��YL����88���>�_2z�$�����Vʳd�ê��)��]�!���*��������j��
�g�\��\u�xiU+��g(
�N ����@�Q�0���Є��#�q��K�<�"�<h?�~�Y.�w��K�~ՊC�����#��]���E}dDĥ*�8�����'���������l��X������SWX�("d�W�Տ�>���k�����([>�O�H�jЄj��ScS}�zB>�.k$�m����z�(����H��D����Z�sL�}c�[�cY.kՊ��G�re���U�d�+i�{�
/5	�<�_Q�������3�0�U� E�|��`�n�*�2 j��:�蜩�f��ی�&��v>~�ıR�m��|%�T�M����Z���4S���o���^�WW��I��{�� �/?��<`i�\�(C,L�����8i75��__�֪'Z�x_b����9lo�ua����̪�+XC7��/��lI�\� �WX�~�j7����`n�����Rr	�b2D�}���P�/��W���(�ۼBРHK�V{�9'=��L��/�TU��=��7v#@�_�hf�k^D�ed?�r8k)����U*��Ր.-G�j'	'�خi�+���*��.:���F��MZQ�������F0g(��d� �7�a�2߃Ez���_�ك�b=��MM`<��``0�Lc�W�`]@'H�/�,�� I��%��P2�dl���S�4+Kae7T�`b�i��X^R�|� a�vc���.�������$7�J��%�_&7O�<��sM���\Ԟ����	�
�@��-#I*��zY�}S��l��Z[�[�ZL�>��Ʃ�1U3B7W�dsEDuc�D:�ު��k\L̒�ֵk{Ym���`#��wi�d_��3���n]���?5�����W:��B���������>�����jD�K�-6՛37�.τci�/.��w!P<���<��||x\�#s�������?��=w��`'w�mj�������[JM��m�'/o%�3��p<7d��P;0�f/q����v��2��尳�c��G��o��X�L���G'~1��K�<(BO?��vsXŊ,���E�SΦ��M9[���k1au�*����8k�9�X�������(AϚ��3��_�9���]�s	O'��3W��
�����:b)[�l� ��Xv��6��Es=�[(^5����� ��&�֒RF�*�_=^+�#�y��N*�TM-�v��;�a��r6n7Kp��jIŲ��GN�X�e|y�h>3����o�Q+�.�}N;�2
$�J��" z�k�O	��5��K�ô{z:r½@��N~��F]3G�#&$��.�Dӈ��ݑ�
�����ƺ<R������8������7�F�]6��]��M���:������ЖN�y�&�i��ހ���r�w�.U�ށ������3`<�\���`Em���Yա��Q��.��v��6�NA��? ����i��{�|#O?˙�fD&��8V����xA�ud{�: �rƓ�V�I�֦I+�wxc��'J�C�j$1S�A-1�\E^>#�5C�k�=j�]6���\
Q^ y���]��<^6Z��W��RcP��%�8�rZ��츑�
�oF��S�������	<eb��.^A}`�U)QA�A���K�GA�p�T�R< \�x
�[,_�����2�#A1c{I�m��X���b�[��(�ڟ:?-��4�O���[i0�AN��#�@Dnf�PH��&nH%�o ʈ�"���?���3�w��o^~��a7o�e+HK�����5j2Dy(����D��=d�����=�ٍi��sm���\��w\����ƾ�e�e�6�(N�_�	�%�U����p�F���� �cc��5}i�W1t���������i{�:��N/�\�|�r;�U�Ѽ�Q4| ��>S�D�6�e1�Y҅��VE�E4�џQ,;��)�Z�&�|8z�A�f���d�s�>�R�%��Ⱦ&�饏�_N���7��o����wFbc���&)���:���x�|��ŗ�����M5K�ԏǧ_ �G�Q��y�K�<E@c?���d�!�A����O!z&�l�y7�<�.0���Ib��k26jAf"o��+�A	@�KF��}c�!�h�w�$u
ȹs5�	�Tˏ�Z>��� j0e��<����>�)���~�'b�K,|r��G		Mu� �����w��&��.qe.r��[����=���G�ձ��x�и���O;7������(_in0G	#�N���`>P���|��!t�B��׃6���]r8���]��KJ�|ME��%��C�K }>�_��j$w��\��<��v����-�n���)�Hd�Ĉ\�OW2���M�\�3fi��]���I����	�w*y��<Ԧ������Y)��?4��U6�(�y�i����GN����Ͳ"�?2T��y�%�fYME��f�|��h�tL{4��U��&./��+l��,0�Q�F��[�����P�Q�9I;���e<a�G0H�H�m�2w�K�CkG.m�v���58<<�~w���'}��%���7�ak��G?��X����WU�+�?��,�E�M.%�Sq��X�����꩛P�D7����a�`�)�^"�Ѫg���`��y�)�ҲH���?���8�P�s�����T?k�$���5j�%Χ��2^�W�w����hC����ZY�b��\�t��Z�h��
�n'�v��5=�3D�UtUAՏG�{S�X2�F
�+7b2�����M���%
��B�[i�];C��/�8�<��6�+�Z�g�<��o�$dd�&;V[g�$�!�f��wt������mY
1F�wEOb0��'?I�N���-`u�g������Eq!�f�r���X��!�51�BK�U�X�a>�x!�k�I�)ٖ�����z�l���C�َ`��Ñ ���I9{�-;o��d*W�m�z�mx��P˯QGid�Էr� 9ǂ_�!g:[��W��G6?�~�:j�b��/=8ȝ��%�tjE�mޛ�m��]�w�"�s���p@�R�?�<#TPC�v~�q�J���4����W�y��{�Ll�Q*�#�������Z-<��<1(���%�5Fn: LE�^{������H����K\+��W������i�ϊ��I�??Ɉ&8�i?�%Ղ�/�$�2z�d�*U�����`�9�ԣ�W��m�ܔ^���e�t����\~xO��f�@)�����0�s�g���֍CfG��]ZS�x�:����lJ��@󱱥K,���1K)���-�������'tj��,G1Y�ڡg�
9N���K$�~�u�Kh�U���|�����9��A3T�h\��\��9�X��a�X��(Y��l�'j��0#��I/ڙ��~�#
�2�>�z�4�������a9'�����J%E�]a�h*�^�\��ԩ��q��賭B#z_��\^5N���F��E���]{N��d�t��N��ݿy���h�ZW��-]����g�.h0�ϊ��r��_�ӝ���D3ҋ�$���	�N�u0���[C
��V�;��Kƿ׆�
D�H�E��'m�+�='Js����z	c���Zu��$��^��-�7���k�99�X���,C�iR��Z��h^��.IȡC�Z�z5��ZW r�޳=�o,�s�7-��s���t�Mb
���9xQu��+�w7Q$z�b*��4����EJu�L$[��[Q�%Q���W�/ZX��~͇��G�O֏gnJ]�m���)ʥ�2/����3�y4�O� ���S}?H�т@�Mxu��fc߅�l�GV���`�|�[f���,Xt���`��c�3tC=�?1�q&b��eg�5l����	xNd-�[���j�u,8�x �4p����{��R���4�퇹�g��Vj��:����8�/I�vbˤ+����θg�Cr�~a�e�Y�6�=&V��D����y�oX��8ʔ߆��{EY�.���g������|W|�! /��0m{ y�$�|�*�(�P���������Mly�	�/Jf~�<]�[�����K{�d�CL�3�6�:tzk�ݘ3�{��(�D��8�2�D�#ܦlV.8.f0H(�lYBB��^U��n��|F��;+Ŭ�1�ȇa����7�)�׈k�0��l����ސ���njyL�Ц/g�Q��
�K�j����㟣�@�@Bˑ�o|B�*0~KI��-�^�V�k��sd���@��������@;F���Kh/��=�����>'6��s��G���@.���K;[[SCx)ד(�\���E/i�'����;߿+��O�-@S�$P�O������_�w&�S�J�c��R�2
+ |�5K�������r�6\ZK�"�~�����*����d�u���ʹ�Kl���"_o�hIŃ{������}rbT1�e?�-Qm�T���^JJ7w!�w��G���q������v6y#,&��W�����np3R�I���q���r�ƣ�S�c�YhT��a�8�K`�F�~�R��ㅓ9�D��!M�Ȩ�?)z _��5�/N�=�3b�������U�cB�vݰ�$��?�[�։�G������q$M�\b�m
[���2�X�Cr�-���s��2"��T�E�=ar>nsK�a�K�?��?p�y�_����>�u�m��F�>��)	W���_T��O��d9������B�Er��o�ĕ��J�K�.���~�~&i�F*$/�9DTQ�wqҼ�\�:e�"��Y�?�}�କě*���3�j�~� 
y���J�L累1�VQ�V���Z@��dP;[ƻ:���(���u��%�/�EC�B�n`D� =8����ር�	�}�t�s����4 sr1�M���Ue�t���'Y)�D/�kke>Ea�$f�1�9�t�U�36���)��I��&;���q����@��Kp�I�ٜK*��hc���B��[�+�4 &��]X@5���,<;(<;W��\�!'��uz�D���ê<���d�%��M��٠˹��O\h����-)`�X5�c��(���}%�yW8��w�[�~�yn���$��y�5��S��Կ]V���O��� ,[z�P�j����{}���x���A��eGW ��A��ӭ���~i�I�|<�-E$�O�pw$6U�м>?�T��mG5Xy
�)++������Hm�P�Nw��ZB�v�1��|@�l�R�Q��=,�R>q�r�I�k��~%�lj>�5	'|m�q���c�+���1@8>�{#Q����*��E�n<.p��K��X��h%���fb�\N����T�e����v@P�w���J#���\C�C_����fmx8-��:=�b�����Nh��*R��rU��k/v�����V�g�j��:����.�$��I/)v�F)�TNW��i���O��P�/ ���D=w�)��>::'ɟ����� ����b��]���н�� ��[��l����3N�pO����H����X��ߝ���tը�MKo&���z7�-�³�P�����7�r�ş�PufNI)�}��������f���d٪/�NCϗw%!��b�����Q˷�-��~�/��������޶���輟^0�д�o�6X{�{��aR1$��]�ǡ��������s��ٸ%�2�mvW�ɓ���`�sW���=�K*�൳�W��h���aي��!��&�������M�g�a��	����v8���L@ ����Fbs���x`>��Ee �`B�ke!P�����<'
��1�A�O��(Op��C��TCb�k���)t�)��vYߴO1��:U��s�;�vk�����	�����ǐ\`*�|<>r1㰤$n��zl�2 �1��
�zr��Z n�x(9�H��M5G����f$uC���������C�p] ��s��h>�ok~ջ��p��:�_.�$30¡�J����1~����ou��;1�F���B�N}�,�f\����}�	z�	�BscM��f&Ng��N��6����#�� :�ow�.�|����G+<����3 ���,�K�?>m�$���p
ic�Esj��@��˳E/T3@���s�T�#�Y;'�f
M���-�lm�\�C�(%�1c=���~�oMev�/����!G��� N��#�j!jC5�A�$aJ��X S���=��:![Eʢ<s?J)_B��(�r`W�[u�/�ůK,D�G������\zc���0|^�F�j�W�&���Yˌ`j+���q�/Zb��ժ����o��t��[�-�F��?�(L+�yB�o�����wy���?͸O��M�}�3�(fsT�v���|�W��2kQ���Fv�����X;�+���*3a��CB�4�,HC|��q8~�J��9Y5�$	
nӿM������]�����44����PV�T�{a���Ǯ��562�o�W��U��.Q�r�,�<�����p�0���o����t2�k½*�A.V&H�dR��"�+46?P2�|���:������8Vh:�^�g3F�:������6Z��R��e���v��@�����vo��ޝ���������D��y���B��5�kk�7�>��3����vӣ��t��a�`ԉ�#����1+��dc[���<�����|�.��r�z�Z�d5�V�4�~���z���H>�RY�K��������[���nn�"���&t$�l�x7��?���6�J6C�f;x�M|�R�{��6a�@x�o�iê��c���l7̚;~�
�>��E��E����.?�@2��(�N�B;禧÷wzT�����ƭ�����FGx��b�����p���4�coazi�{��H5��D-�D��XE��@���ea���ַ�O�����"�����k��ǯ��:MJ�m�C�҆��z�t��ɭ�@[t��/t���Z�����&�]��LK�m���������d��R���anGHr�p�PzaU�����6 �d����/�ߵ��9���`z �m�1W�ED�8�a.�ȿ0�
ݴ4�=0��<U�9_R�#�������$�G0a#���}/�W��Tx^";��əߩm�jZ����E��o,]^Yb��(�GFc&:\�bi�K�w��������ݻ�K[Z��hB�9��I�������k�������%u?��/REB���d�b`X7�����˂ڔ��nǗn�
�ښF��f��?-f�[��@�n�~M /o?���1�Ac���qD� ,lKߴ�6���bD�`4�Y���s��Y��*�p����ԙ�Սu�yky��!'u�s�3����|N���ك�/b�C�f\�R�J���D��"�4q���7���>��L3 ~'��O��qm��Xǉ��'TyS���l*��I����z�&f�i�C��y�Z�EM�_����/P|��o=5\}���}�?�������ts��� Fքa�_dU�[X��`�{E�%x^h�H���5D���p*��kǚ�I�E_ء`���-��I��--�d����<V<V����9�M �J��뷛�lU��U��I��Ĳ��;��X:�k�T�t�Ay�
<K&.���ɾ��]"Ji��������kM�qp|㿑�a 
,OK�A���o�*e[Q8)��jg*8q��R�ьI��?�f�WR�����銳�䳌+���f��~��_�.(�%≑Z�٥��(����~��%&] �R3�J��Aд��I���l�Лh�E�O�+�r��X�&}v4�����́39 �:\,���Z-��>%	���U�`�T2�J�y}}��Ј��PK�Ҟ����vu�8K�\��S�]�����\<�,'��]b�<���㈄ñ�]b���s�z�&ޑʘ7p�^E�u����L~��=�� Yn���X��5�j�U����Luv�S���9.C.RQ�
x��x:��X��N�=���j�A�����lQ�W�?A��Q�N�8߲D��/�������6�!�n�j�d���V�N��h%oIۺ�>> �s�5%u� ��i��L���5�J\��T\�A����a�Z.u�Z�������k%3��,���xE=*��D�Ù�]�k0�F���-�W�p��A[��M���0��'-��������
ާ��B�7L_�#���|4�hB�$�K���2g�X>�������H�$絝8pl�!�x7ziW*��LUٌ� 6��n�E8�k�@�uC�.��}v!I��@���9��µ���w�$B�2"�Jw�o���"�������"�M��,�p���u_��H�QˑZƃ�H��2*Peb>��B!���J پ�svJ�>��q���}6^.�_z׿�n�IY�/���m	��U`�A '���	���yy3����3{�v�D^�T��@�y�� %L�ɎQ(ƭ�����-�~~�G��ag_��^wb��ZU�!τ�-�u츴JW:�췎+��@:n&Y�@��o��Ѓ��kF}#�o� �i'|����	@�V��8@���_.��[oe�4u-ݙ���X��%�輺6J8�Ʉ�v���#�?:�N�����P����fY[�ψ�dWY��Š�U� =I�5�t�o�[��v�o�7���4��K��h���q�dQ��F�G���U���U	��zg;��4�g��/o����5ʘ������L�M��$�:X�Ɇ�[ԳS*{�7�	�����d~D`į��a�77�"q�d�0��{v����g�UU�F��4!&Ą-������7*�+�77�w�6����bd��~��Y��MbI��`,���N ��v2b�����V���+]�`�6���8b1t��R2��'*b8��O�*��7G\r>�?�4�?Te?A��d�ʔ��
��F�j���M��	��%������￟��@�]�ڊ)ǋ���zn�Ɣ�J2���ӕ���/T��r�+�"���P:n�`���mﴍ᳴�<+�WT�R!��*��?���>w/� ��7xZ������qk3�+� �A�H,��� B'�L>�t*��+P ş��"�+�Զ��E5�E��S#�0��f����
�ê,�\}01`I-��T]���;�^?b��	���O���;B�*��+u���ZBSck� A�g*R�ϗ����N73����j�C`�C~̯�g"	,�O�X��֣���F�ʏ�����Ԩ��?#��pV}�Ow7nP5��wIP� ��4~���:�����*JUP5"�F4��# ��8��ΜA�&��y�!Ƨ����&�wY�gZ?��2ө��ߩ񛂀���N�t0��o���:x������_��hV2k�H'wz.����Gf�wҠ�f�"��H�=i|�(�q*����yX�	���+	�u�Oa@[��� ��6���g�1�=��:�sL$v�UO��<aŰ	�I(I��%/����x��>GZ;e0(q�#Р=�λax1и ���"�4���#^,!�
fs^(��I�I�TQ+��n�t�-�Z{�ĵ?�3�@o�� ��$�E��H�1�{Q�,�@`e�3���0$��u��&������Kȏ^+\f�<㝢a�4f���i����Y}����Ʋ_`�������*������x��$��3�r�U�X��ߝ�""���L��_b �8�PҎg��^M���&iB��8�,G� ޏSu�ȗ���<XSd�V��u��
*VJ$���*��ڥ_�F�9=�H*���������ͥ�Q��1�Cg�v�P���uP����V�/��<�M�	 f�4�}��ߦD�g-��aq�o�gCr6wg�ިB,�v5?����^�C��"kG�u��jXkæ���M��uJǇ�����)a5�en^�(*]�\^�2�/���  Y��yX�] '���9v��nP���6��lc���!D1��E���p�-�ȹ0�b�g��:qs.u,^̦��>��F�tߊ��Rd �\&0�a��律]�;�!" ���KF>�]w���E٘�:~�i�fX^�T]�F\����DY@��� O���w8E2:��샽�X`x�`�c�hm������@
��� �]��2?o��UPÐ��2DEC@7��3k�m���mL�K�r���~e�ټ!�³��ֳ�ĳ��3����U%jd��sur6�{�B��%�L�_.7u��Vg�lp�߿G�`����2�g#��7޷�n8_D_\½ �W+�2V}sD�pVK)�u��qm5?�B&��oa`����� S0����8X�E>�vT�[B���K����6{qwzΑ=X�_��6�*�&��X,ݱ��3F����~��ҩ[x��-�Z_��S�X���#9I�z�ѣ^���o��߼�  �~�G��1���O�[�_�:_�n�p� �9������#f�C�|�@�I���v�Z*MQ��J�A����	v���g�{�_%�gh� ��]��O�|�ȹ�������_a��sp_ +`��q�b�q@���|�%��}�P%d7�"�4�	�������.$�l0����z��+�[����TR�.Mmߢ�Fb۲�Ӿ&�Q��7��� ��������e��%8�&��'�X��Ey���A"��o2asꗱ���u��dq2�<A�d�5�9y[W���չY�u��P��� hYƘ�L��I�yWk�F���:C�3�LRPe0��݇\؟��+�2|FL.͂�,/��J9_S��Ru<��D��F>]����G�ă����u��H@���׎H(J%2>���e���ؕ˶��oWy��[[�������:�����	3F����}:Z���n�X}��'����RMKٞt�t��U� e2���b�᳛_I���[�&�-��57;����[���X8�S3��v���71r����׏U\���dx#̽��T���)�M^O�N���oᙦ����tR&��E�,㖕�m}AŸ����۷VF:`�#�ޓE:��b|������K�eJu{e�2��;z���嬃�	-)%�F��ز��$���q��&;�ψ�%r��H���d�f(_�2�B"�8�u��/yϗd���� ,��̌Y�!�{�Z���Y(V�i���_�&H�������H�e�(�"BK����?�mMx��/|�}�M�#��Í�:p&]�bG��
�}��3�2K" �#'�mgm<,V�KKdv�>�=j+H'SJ��J��E\K�>�s�����x3'��������G���Ã�
o�5B�m����B0�dKW�u;��:��E|`b�|��a��D�*�Hjh�9��������vg77��>t0�E�&Ȳ�,�s���䂏K�����L����y� �����D)p.���B�k#���/�o��W����O�	_�j;�h��o��H�]U�MZ�3h�9�~�7K3�3 (R��U����<�ckc#��Z=��-��S��8��l?zs�_���n;=��O��z��w� E[��i��k�t�j,��9z�CA��ח�Eg�h4�宇Ҵ���ԘwU���>yT���^q�����5����`8�k`�r��}Tt���<IT�C���[sx-g/��FN5�e1Ɔ����J���� ��G��7L�B��;E_�s�I|��>���v4�3'��ܰiz1�:����r�P�EN~L�=	�i_7�����L0�Ot�`SzO<��T$�:SK�GZ�ۏ����z�8a��w���s��q�!}��c\��Z>��	�<ٝ�mc!p�E�<"/�(�*���A*��ƺ����_�-�%-�Vj��!���ӓ��i]�ؒ六s����u]ar�⛫x���˫��DPP�t6P�1;��WsLz����\x�~�ȥ���Dk�k���Y*ƈ��4gJ��	+vO�ڤvtaa18z?��e����6ƛԴ�O�8����'S�'Sm�o����d��BL�f���W�����@%xR�����uAJ�����}�WC�X?9����%=�Yq���r{�ZøQ2�����K�V��D/ND\z��be�8(	�ޜ���s�+�g�j��"(���Y\��1MR.��$*kK�R��|��\�P'6�Ƣ�l+}X`�G�:I�%k����M�$�d����G��YL�/ON*V(!�����u(��o'HX���8��_;�@�b�OY2M�A�8��uy���T�%����HI1�j�%����6�F�P?��m7�L���hr�>)�Llmv
�?���]�����f�M�KQ}�3���`�孌���$��,�V�G>#�Щ���5��H+���
�: ?�wwjI�J����C9�k���;�CM�j!gq5�/ȯyC�
��uJ@�ܱ��@�\�L`���e�7 �,�����$���6*T��仴�!>T�r'��A�s\���P�y,g��ĳ� PBmm-��S�ti��	+k��'�vzPZ1��<l�E;�P��'u�Q�O������힕T���7�E�P��N��,���ٹ���ڌ"��ؔz7�I���xG,]�:Ы
�ۧ��]�P����QK���ߝ�Q�;[�6��5�_Ci+���vk�����ۿG��6���y|v8�x�|'��Ϯ��>I2>�=�l?�y|���;qC>j}������^��k[�������G/?>-��.t�����ڸ񀜘����؍|9�"��D��Kr�����b�i&s�����R���l0����ݦ �ͦ�}��ur��$���ݷMخѧ}�x�����{����͠[b�K�#` ���K��Z���&�O��L��屰�ș��hG�&�V� 857G5h���|�:r�?��2<,��'n�Nx�C��^�縤|8/A����L�9����(ީ�耀.�2(}o�9�v�-2�A���0�]uyES*��o��Ь`�b�ʺ��b��@O�v�LT�D�p�F1T�=Rn���Vt�� ����p��:�# /T�o���}|үg7�����j=�3����I�UM֠�M�[��.�dp��m���3]�B��'[�7�����z$e�_��OKW),�	�
F�	�-��_o�y�o���⻠-ԍ���n��<A��(���:�NR���`�H�_GC�g�л��;^r�����9/�&v^J]}SwA�Wd����8��-�?�$0���}U�)K�{yƛ�����X�Ъ���R5��y$r2�u�r��û��\���S�>�rh�gs�����};J�{�^���ż��L��qw�N
EmB��0��n�KF��r����z^&�4����lTRI/���#\�P�����y���yyy�M�ʔ�t8�춉�"�� ��II��L$g9t"h߮���]
����w���70E�¾h�ɦ>A��-6wm�'#�Φ�Ni.�5(��r�=�������%|�to
��ޭ���S�����5�a����[Ȝ��BNN�;��:����!C�i>w���ȏG��W^���2�747I�A� �$�~�v�;��hͥgTO�C;�4�g%Y���z��G<��
�Qǽ�� D�w��N����$�.�M��f��N0�
	��h�F>���]�L�P6�V+��C�L��P(�ɸt���P4aɯ-���w#�V;�>���J��б8>kMl^9�Zz�_��5����.�~R���>�K[��7*,�G:4ǣos[�jʫ!���X8��m��ťY�|� <�*6O@�
X"�� iVYE���vF���c<&ƪO���󑧛��,�Tx��+�6I��T
8�)L�Є۬1����D�S���噉!_0�	��P Ñy�ɀk�� )��������Ic�	ʮ|������v�[:�>�����t�B���*���q���?��+���r^�5���P
Tr�"!4�|޶����O�7��[y����Ο�ܒ�$�x� Y�{&��<}�Y�w\a�Q�sw�@���n�:�QeeSRX�f<���죥s�c��t�[��x}IL�zR&T���d%%�Ve��#BN5�P���)������/_\����/��ݿ�AjF��t�r���t ��L+�}���wplE���lfJ^6�#M��t?����]N�@�L*a�R-tBq����z���?&�[/�v)/�^��Y#�k�@ۉ�ȹ:�D�b3�Ǡ �xx>̉�y�0x
B���9��LH��'G�jGS�tk���ֈ�t�C��u��`���sѱ�̷6c8��c��{���}�!��ܜT�OPm{���=3 G��Mկ{ef�wV�f�n�-��#��������8���%��m�Ϊs�$9�=��2F\�@큔��ӎ���r��B��-�YK�O�^GJͶG�FRk$Ԍ1ӕ�l��N�;'t����ǹt��|]�p�<�::����4�U����wv�Q�Ƒq��fV�������fp�.����X=(�ccY9h)_9�yt2�^��%�6D7!�K�U�*`T�λ~\�0O�]�T�voeyX�'��z�z��f�t����K6�Gېs�J��
?��+����m,s�wZ���S:��{W�O5
c ��VU_^�5��mw�ꌋk�2��m�������޾��>�;ۉ�|?���ANR;|޾�+�.�q�}�yϷ�	s�$p�����-*�K,߾��8�D�K�#���u�u�a7a���0ziw(����{M%�%���(��x�N��L4�f��~�ڧS_�K����֡�Ӄ�'~!K:/�1#5	U�K���BO7��vvU	E�Q�v͗O���[ӡ�P���������L��ݓ��;��sǩsǧ����R����ϛj�Y�R�I�~iF)<�S�%|�[-??�0&�At@���dm��"9נ����G�(֭2�ڵ9g�ͣկbi�>�!bS��6)\Ȑ��@
+/���:p�ڥ��8z��*��9�x�6��i����T��!�G�@[�����/���>��=ô�����yUҢV�/������ V ] �Kj7�5WU��X&x~�L=�����L��#Mx����)[!�fM+�o^U7%s�`�{;���|��ؘ	o�%��K@���;ۻ��y���p�~_�����q�;�͕�� ��K�VU�����"���D1o�r���FX�ƛ�r8��; Y������#_1���.2����K_@p/$E�����n��&i�V[p"70����[������#��/I�Ǧ���r!��㔿��Sm`o��1yba���X7ȧ,�l�TN��e,�u
�a���^����J��=�h��3�`'+�5j�)��������S~��Q%��>�{�^����f��#?&�ck�ʼ
d������ԙ�㕭Q�!>.����_oo�V��l ��Mi������^������>#Զ��^��@oO�f�ϝmN��	����h���!D#���	,�,Lt%$F��ް�p�Oչ�zU���.��jiU�������e5�s� /?#^;�����2_E��ñ k���;�e�����I����*z yqq�1�^�坆�e�僋,?�`>o67��mr��׆4?���ؐ͜�;w�������r�tR
���eo���j��\�[����s 9��f FP����1X���v(`�)\�LaW�z�(�D|�#�^_x<��O$�̱\(�'	F����A�����ll�G'a�y2ds�͏����|�(�٦���P��,�Mއy�ϯ�l�f��!�����q�k!���0����⑭<��F4!|��2���qC
#����zA>�ח��ה����~Cl��N�!���]��݈{��.6�Z��eSQ�e�C"G�h6�O���w��8z�
g��?(���`L�&q[gٹ9z.ׄ�֥�:/i�㘨wt�bqw��J��P[������CF�$r}�o�\�Khc$��P��<�u�nbl�;�6��q�2a��&�����F�oٯqJ�q�ھor�]���
����9֪���!�w�U�j���G���BWN([��"��i���j�{ꔃ�s0Dn�.�O���5�Um��_�D�������E��5�Gű���H��O�vz�ܨ:x𢨳��zT5j9�O����ι��t�4�$� {W���xM����q^;~�a���\:o�O�_O��.\��������_L9R�?j͙a~�<,����v��>����刾�q�һ(��Pih�3]�Ү��k��sr�r�C��ǯq��D9D�|.�7���YET�7h(�P��	��ϳ�EhR^EV&I�3��*���U��+�Z.���3��$8�����M�Z�\9��d!!�d�#�(:��A�ĉv ��	y��ıoԯ����һ�Q�vo`z�� S��Ҫ�`RT��5�n�5����3�|�j���v4K�/�����z�7���F�������,����p!�||_�RC�Qz���8��l�5�0|׿|�OF��W���߈�R�+����#�{�͟Th���vVG�U��@9b��?��c����-	
�S<�)ҕ`��G1��K��~�8(߇���_P�kkA�pD�`��A}{;{��[[�����Qgţ5�!��:组�A�_�t_���-�P���f�u�G�%�^����kt���BMj�2�O���3��qK���`�n����:��q_dp1���[lm����7Z���=
���j�̶ge�,�����d~?9�w8������R^8`c/D5x����D)󢐄)ތR����$�}��)����@`i�����@+	+w��qBH�3����Y٪ै'���_I ���~�s����0x"��Ҕ����������o���g��8�^/��%��������yԭQI�H�|�M~�����;�7��B���_�Ƶm����\O�����Q�Jy�*��^�Z�	�ْ��!�����'��ǌ:Bۻ�gp`HӃf���V؇@� _򽮰N�T`��G��:%V�go"7p?��601����r��Pi�%[�U�m% B��,U���ee����b�cV�Ֆ�����Ӹ���-�v�	���{�������r�;h�.gv5�	���r�X��4x���Fw"���W2�e�~��Zj�����Ì/��c�H�c{@�Q�P���R;��V�fFb`�Vѽo�RO��[�]N��� mCG��E��J�#c�&����HA�b��ț	�WU�����u>L#�k���`a��"�t���1���
u��6Q�)��ݏ�q�����`k]n4�ISe����7��i�S��눕����u`��N�3���¡}�n�҂{�=��#��T�ȭ�om�bh��tb�7��������pr�#�ǧ�֐(�.�&O�'��1>�&�/��Z5 p�B#��W�Yµ"�ƞw/	��}s�����J�^=�=P�9���c��S=$~��s�MU�&��J.-�汧�R��/>�Yj�D���.猟ˌ�/��+Ǟ6:C���]�|,��ٗ�/э<+�����3��Wk��������6�]7�N�kz�>����.�G�D���C0=�u������6�����:��Y/������Rjz�(J<LgU����>��Vʮ_"��&�(�!�(Η���=\�ͦ奐��A���H�T×
��^��(��`X#���`�����ތ=e��D*^KE`s�m縐@QU�*�9RQU]�{Eޜ��w�;���Ka�[�FKW�������#%��w
Bkb�,yU���+��>�����y�|�i!U�!��k;���Y�f��xi����L�'�p��śu��/&�R���1��R�ڕ���h�gR<9Ï�H	���]=�|��
f��x�p�L#j��?�Vb��cQ�%�Dn@�PXG��j�#;R䪨��+�&2d�nA���m7׺o����m-&���S[!y��)�����ɠ�Y��4�G�&��8�/�z�r��.=C��ag����=|�ܨl�3������!�3���	���Y;OGRA%��J"���P&_U��+NP�����;2
��E�.�7:ᨹ�}�u�#PM�n\�>��-ܽ�1/(,��p���&�Pgs��~	G�>���ZQM��&�h� �/�ac�����6��7��Y�l�&�-t���U�v��ŭ�����%��~����ݿ���I q�o��=7j��5���d��r)��Α��s��dn^�u�c�� " ���6��yVn{��+h�&5�Y�ge�J�����
RL" N���f��C��KK08��UTV�2���X�g�;-���5�הL��;�>�Iw3���9��v��& ��j�9Q)����2�ʘ��p>��)ʱ>M�v.w����h�A�Uܛ�٪��U������������{]!�mx��z�O2m�O�`�3�k����`��y���bPm��dR��̆�i9{�ˋ�t�ҟ�����@{����&�l��:�'��ro~b�*�g<B����?� ����*&	�P�L��ftz�$��5%���ĊH4n�c�;X[�\<hԿ�q�\z��z!��;D��Z�R@8oj
��;�A�;`�q}	�����De�M�g�K�.ǅ�&׎�g�K7Ym��h��@�n��06��wEq���)P���:<u[D�21tn��`kʮ���e�~�2��̇�4	
Ln��|��9_�'�FJ��\�[�s�����N�z=l-�I���^�H!��nboЛ^̻Y�Tr�]Ü��໑��ϓ!�Ǫ��3��=�Q�1�(��vq���׾�X����k�K��z�W�̕�!��P4����dcc�F��L�	������[���,b*?:���-���&�Φ')F���ke���Ѫm#�d<���X�6���/���u���kj�'���S��H�u^~���<S�% ���F���NàD�U�����"
�X_V��j(�9��G]W��D,�𹠗�vѮ�\���y�/�1�K#�C5�Y�U�-��F�W�+��2���_����:bօm�Z��:�Y�q
`�Q>��exPPӤ��y��q��9�������F`;a6�>LNX�~yB�C
-��}=�]5jiP(׀S2"�b!(hds�e*���>'|{΀����M&�x��r������6*@$��v�cs����I^'f��	�]�"!mK��颒�9�P�/����g�sgp�l���e�w2�v��]�#���Q5�!$�5f5������3U�K�}�������Pj�Q� ��e �Los0���k{����Y軁ڊ�2J�\�m�S��b���w �;T������0��-��q��Q��{�0;�n�8��w��4���!پA�Crw��%���
���@���}^��cϚd�����IK���v��.�NOK�,]JRRX��oy>��W�|J�8^��3�NH��(��E��KXk���:O���j(G�Φ+X�>��ab9wn��ĵ����nTp�5��P^��g�JĿ�97м!���Ƈ�v���G�]�w
d��O}E�Y�#�7�=�<����a�%c�DB�N���N�z3@q<~J���\�qYҏg��{D��6Շm�m�=O3F~KJW�K�e�S�7	ץڏ�+������Sŗs��|��%,�{��i�y(ť�,G5�+�����ӡ&����ٱ1����UGV�2e;��H�Z�*J���1p���X�ӎp$_�ͮ�E�og�\�1�G�U�w fݳ"T���o�loZ�©���.J���b|'����(�,�i.^�o������Y����/��4D��&�W��*Q�68��R0�l#����d�_��#�c=�R�P�>P�e�D)�`q�0����633_j�ꯡXy��%�y4c�@ϝ)�mu)�ǩ�z4��ς73�j�����l �n��cJ/�2�A(cHߐ%&����9�=Fb~a��dIF:))��2A+�0`��h�|&*w���:ufyYT�/�����0��$��?���#��1����WZ�,^I>#+�">�Me}J���0���Ua�����޻{�	��ā�>s����}Ƅe��H��ڄ�/�`VZi�?����@�",໸of�~Dh�x�QCH�@w���U�"��V�1�yR�"C��'ҹ�H�S�1� ƨz�Z�Vd��ƕ
pݔ֟�/�@5��_�o�U%ʹWՔ���>y�҈��1�O��2Q��47? �"��o�j �͸�f5l̴�R�o`Eli^k�BA�햞�OL��&��9=.��5(1AW���n��N�ێ����͐�gZ>ֲ�i�cM^U�/d9n�z�[�1�k^�ஓ�}�ۆ�t�e�w�����8��(nf�|��9$c�c�߮0>��q�������=�?�_/T��hV{�1!��/W�ZLV�u<�=���K��Wed�V$ �2��[�c����;et���.\�����٬�հb�b��धl$�B��H�>q�C�'X��2<	��;(a�r�\[�_޾Śv<�w�H���~����|�bk����QM+r��[�c(�^��_����r��e�<$Z�3Q}��(N�2!�M(/����`*��(n��=^j��l�*gx*�s��H83u���� �!C��%u�b($Z2p�)����m�Sej0�J-���qt��L�wF�\br�[�Ć�Cs)s�uC�-��~��KL�%1��
�����%���Q�ro�~���}{�������|~����\��ia��NhmUp��4�[=畢vzE�ǌ�en ��Y���J����0�Oә��6�S��h���옎.mˇ�c~O�J�^r��p�y )��w&�Y{��X��I���MY�z!Ea)dQ1����Q)P~���s$�N�g�V��xB�s]_��VXeA���B
շ;������eskq ��`΁J+z\���vĞ6�sz�������Pe�NQ
������%��}�GE�F}�]ܽ�k���aϭ_QL��b�)/�&=���F����Ú�OFo	��E��a��/<z=LI�W�/-_�.��.+�3���3h���T���o��￾<Y3'F���]�YJ��qj��m��aq�9cN��jA;�z�����q)VI�g9���`u�����1{�,���7�~��i��g>���j�}:6��SD7Stf�����7%PR�����mJ����g#}Ȭ�D��b�g�h?U���۫�&t�b��)�"#nϡ�C�A���>�Ł�*��x�޲:;
�uW�pw;Q�j�15c}�:�)�ksn[FC�/xi�B*�M���R��XP\��C�������ئ�n��3�F��Ռ���l����љX3�Jٹ��WJ�i�q�E�Bߥpo���|������]\�g���g|Ј�ц�������,8�1�����'�?�^\���t�����F/��9�$�߁(+Q�G�PI�j�we+B���l�dIYV�DS�,��jX�����S�5Y9Vu�Y����Y��������N'�&<� �4|Xh���#�Ǣ�fЯ����AqN���
F��5TW�a��|l�=4�Q���4���"��h�d�4��]�T)8pN��y��'���$��2���?��Ё��z0�y���1#Ϛ�>��U��-%Y�WO��sn习�_OA瘸� �s"!������=	���-��ܵ  ����K'�,��yw���*����� �f�1�g|������*D��c��x��u�Y?7�r������g����j΂�Aܖ�Dy� �+1z_�}o��������]��~�q�D��",���r���Ǣ�m��&<�~�w폖w��9��\���H]�K�".B�~r�Hm^4r�V�~�0J6�\�O�9鑺yN�n5�k����nu�z�`g_W�	*�M'�}��^VP~)2�T/T�{d�ה��*�6�;bQ����j7��I�Z�@��������E���{}�"5���K�^��6E.��,#j�!z'_�x�[?L�
�o���t"d?�C~m�β��Ğ���
��G¨��
$+`�9UĐ�iX�����Y���c캁B���:���0�g8)Z�'����*w��W"�k���
��:�
PCn���q\�i�{㗠��r�u�D�̛�ճEֳ��@<X[[�H�1��]�h7(�!e9��:td�#p�yS��KaW��Kz��pt.80t3�T��*�cA뱛ß I_Q�N�2�¯�H�������$>Y�m���f�k�*�A�dЖW���W���,_�u[�J摧kh`��b��Ԃ�DNkkoo���т�V�^�;R
�Zy]�NB�(�������wǦ�?|�G�z3��7VB��:Az�4-��'����Zw����ıJ(�r����[�k�~�C??ęT1����n�_{U��nv��t�1j�������v$gMͯ���;J���2����-�ރ��E��_���"�W���A<�-�ɠ�m�%��S�fx$�am�$�O��i��<*��WKF�>ONNVd+���Źq�|v炮	��L���<�Ժ
 ����G'76(��5�?7�5CBm.e.:�~�!��=S�?�G�%��S]�|����*Yj4���&��ٚ��ũ4~�
��٩L`p�)�|�0@�ҍ����o��AUr �BQ��ą?.�/ep@
Rn5�o��8���pw�θ���9��{��ML��'����^I/��ҿ����!��uMe�cc\�li��A������i!��q��k?�k�!½���%#��_��GU��8u��ͤ�f~87�u7���:_g���9 w�0�<w�6An9l~=�z�q����Q����D�=y"���ϝ���zZ���tF�)��v�IOY���TpouJ�T���z@kͶZX�m�M�;�p?#\���	�2�m����Vu��ۉ`�Ѷ�N��V��0j6�_n U�om����S�u�w�˳F#M�?�tK(m�\�>2��ل��f�K<7[Bv�9V�A���x�u跃����#�5r�m�?p�]��v������$#7�`�+�� ����K���ӽ.�C��$�e�����6���#)A��|���L�{)�0$m�Ӵ����N��}$%_*T/S����[�qO��߂��ݚj�������|0vg��h�"��$�T�y?�y�rÞ�?�^e���9��;6{pr�����c=-��Sr�{�V�d��3���2 E��x��qd��B_�חI`j-x�b�5�mt�|�	�B��u	��)j�Gw�-!dZ�c�å5y~�
��}����9-$�����V�a˟���n�
�G�2��hX�57Oڔp��1�.\8�E�u�ZKw�YNKk~{!���Q�^|�OV�Zֶ�5§�c�����vՑm�]]�D0�� ~�=��z��#�j%��Hz��%�~ҧ��p2��V�K���9\��|p��<{���u�<�vj@s"�N��e%V���1�F}��+1��t�=�DV-�����ꝃ����"�6�@d\!��Z5�U
��8��k���6'ig%�?_���!r>����;Z���>��� e̯d���m7���v]돛�T�uGo�H���#G�[��(yܹ;��D&T/��@�u�jW���v�����G%O�{�!�@�H��`r��QP9�d�i��x�]#����I!>��Y����7���]FT��+�x�RyW�Ѧp����V�W�AH�[͈]�̝��n�3�H8@��v���Qo,��#v�������`PH���OKO���Bey)Z���׋J���pfbJ�Mm�J�1�m���!��2ĖΏ�J{�h �tAk�H�̢
o��Z���7�i�y	(?��OG�Td<,bc��V,���8k��msq�h�f�t��9��g�S�Ҳpߪ�ݣA�L3h$q�`?�����GJлv>1��>�#�DQQ�r�����å��K��(��-ϩhB�ͽ�ɣ��ч��u����x'nj<���T\\�j$]穤���v��Uq�+�5�xg:�`����{T-�}��{J�F�(�+�>}����ׯ�D-����`U�F���,�x!,ܾ��xL�xC9z��2"�^�x��T��Yh羓r���qJ��	����4��s�/Y��6�ɼ�ҡ6�p_�\2�����$`�(�U×&�<��B#gۭ��f�hvrl�-����u{5�U����P����:!8��N���V�dy�*�`��ǚ$ds����%f0���[z������
�(��(Q����1�@�Ύ�f��yj�d��G"џc��^�k����^���4�w[=��R�C&w#��%�so�(�m�Zo�x7���m�wG�J+˙�2|&�Z#�얊�d���h��K8�N�G���g�	�غ4��E����ǋ�Ǎ��q��>}�4z��a�w3��	��1��VЧ��G��$^�����K�G5�a+ss���M�ٝ���~ �/K#w��'�����!X�4=R����k�;��CZ�Z���0{�������׻`[~հ	���@�f�nG���m�j��SI/_�L�_�'��#w�ӫy��D�X��ͅ�8�}�A5�N�F[��w������h��|8���2I��)� ��H��UQ�j�w��(����Ŧ#8i��KHJ�`as�GE!w��7n<z��[Tʏ�c?���Ps����3���u��Q$2�,XG;K<X���A�yclo����˩a
RL9ͷ㨪�"\UKMI�8?ksv�Y6}���גI���p梇����H$`�ށC�[qx�ğ�
'����~I�˵�����8���k`�f�߿_�α����	�02@���>�vV~����b�g��<Վҿ�X$\i��pi��}���k���,,�C)1����L�=Y=�������%�U����Md-H�,3����BX�����q[x��ek��&@>�5{�[��~��?���$�[g�~���z�8P�����%��r�,i���w�:.zw�����ዿ�g�_�GGv�6���^m9�ݫ[���\'�@�6Ú��c4�#z�=���h�fȑ�j����V��� ��-q����q#�Z~���ab����I��ڋB���7��W�uB��+e��vDX��u~�3xk�1
tݏ<#e����Kp�y������;LT�qAQ��tK��a$�_~i^w4xl��P�i�  '\�L �Q�W`t�z��9��� ������I���jj �,a�O.x$GFxO+���4��C��;-lUW�cV��=J���l���>�7�����6��to��B/NU���D��S�96�J|?�4ƅ��9C
.�e���ćk��(z�4o܈��������y��|�%�-���l�D�c�+��ܴs�Q�J/N8�c�>��pJ�&�mIE_#����N�y��R9�Z��1o��C��A�kx��&D��h������T_Ot��8�i۞��n��տ����1�3��~H��U�7���$�U��W,�R�k���if���Z�B�%H��W�OQs�<<A
�?���Sg{;����� !��{����ݸ�D�fo��tnP�r���|%����'\;G�.e�}p���
u5����KK�Ńc����r8��C&����D��7U��a��n��JǶVEM�B^M�;~)�9���RdQJ葴��-4�-�&�^C�cqAw���ok�1[�����O上g>��]��`�q-U���*�=�o�Nr�2����Bk�+++��ҷG����n1/,���<�6]���X����x?
u\�L��;���1H�L'TWx���~�^���xF�n�7J��`�o�S�H�*Im��/���m� ��Z��|VF���@��������=�mdG|;i��Y*̶��;Ȟr�n�1k����L����b��f��N�2]�X]>�C"@������Թ_�=��=���<aWΦP���8��
� � �*VhSS�|De����I�J�s�2���	��'���.5#C%�m�`C򫯷��u��J�z�oU��k$�ާ��$[�G_��� �����4~�j���%��1S��e([�fIɏ%i�
�B�
8ӿ@�ytھ���'h�Eg� y\�@���A�\��ǳ�(6����+��(0�� �t,?�?'`�.�fAkn���� ���'����v)�qQ�;`�d\Zд��#N�NJ8ŕ[I��a�<&J�������?r�Z&���7���.���*��:`�%��p�v���Di��	�Z${�<<�,�F]��
��`�|��Fo�2h�+�z���"��4 �=��y�bպ�,�	z=V��4�G��� ×T�&4,�M�=�k��9ބ �/��I�i�"�1%,Og��_��We���$}����D�9ωbm���ۙ�"��ڹ�%�PW��ec��g��$[��P�'�v��xB,�%���,��w�L"�
)�'���;7��FS��:a��IE
�vu oyrΐ���diE}P�c�t�a�o��x$Z�7�iO�yO�a�u�S��z�e��p-�5>ԕ��$d&��[|�kV
*knO����D��%]]B�������j�n�J�~�1�F��:�@(?=��|�Ѩ;:u�#���i�s}WcKD��0[D��D��#�
R (�0篶�j}�p#�Ee`����Sլ�Z�S�}�=5)[�O8EH��/��K��Hz��ߜ?�i�[�8����p�s��+=YR��__����^J���-���O��˶�`#���8�d������w������+���X�������5��'���=R�\��t�N2;G����NH�#
��,��ԓ�F��,$��CR�����'g�DЖ��PJ�'g!%kp������T-_���/-Hܘ�@�8HJ5^B6I2���d=ʵ�̸y���0�/)!�49�}�"��f�E0Z���������=�&�����n�����c�O�P��r�x�u�L�ƶJ"4��
;hbtd�,V��@��U"��WG4���y�yn&n��'ci������T��D2�������[�������ٳ�Q�Wb�
V�C��A�{���R�����H݉~��>�v�����s�tm
F;�uj)���ɮ�Q5�K-*��K��;a5վ�Նi�g�^�L9n:5:�Q�#�;���
[��c�t���m&'���\˽�����G*��xdI��!�X�� ��$.Y���ɢ'���u����ю��vwÀ�z��",?B�*���l�s�@2�ӏ��p"Q�ݖ��]sä����3�3�>���z��@K�S\:��d�U��M@><X��i�� t'u(������A��+mc�<��W^r0������k"��Դ	)�.�R�P ����G]z���ŉ���Ǡ<k�3�@9E
�3d�S���c�_�oҴ?���<@G�>Du,��)
�;��$-�Y�HF:�<��`u����4J���a�����moo����\�	��ɲ&�H��r���b&�]v��oq!qN��	�քw���oC�Xs=��̗xs~���J_�s�6C<� ;SC��$��#��J�/�Y�N�w��\�uTb�@Nͱ�F__u~�4��	:����}��,jv!�m8�6!�#3�m��Cє3�|�Z@�S�S{�����%-�}zC{�qܒ���v(=0���v#e���:�;��G�6h�_��:���Z�31(Ξ]�B�ɴ��/��g�0{�$��zs�Cכ7��k#H0:�e�Я��~�r��|A�Y��=�-%�.���	^�{��v��A~�_?}@٫�>i��!�U��`TF�]�3���s��nd>��F1��E��T'/3����{�Gj�Ժ3 ����ꭥ�� �т�/���]�lOB�V�n�|��Z*���ߦ@\?�yO�Ӵ�~��;����Z��	�n��a6���P|߯>Ӏ��{�\��MG��hۤG���Y�M�2Y�~���D�6pVok���tOly�`�AXfP�p|�FK�Bo_^���A<�L�G$�-1�������8����y$y�"ȵp��T�tPN=�»���b���O���\_��I#Mm_��_}wK4+6�2�l��c�W�i
��ȵ~��0�y�:�����1�H�Y$�燂���̞��:��|u��7}F�{i��!*F�Љ��װh�u�&�0�Ǟ��yc���x���nYj��_�¼���/4��*��n�zrMT�e���_,���.(D�����Z˖��"P�m��c�!=�m�$�1*?��{!���=�W�؝��t<�\L �l[E��}�������>�1�2����C�;��iۙZۆ����>n�o3�8��9 $�h��7P�(/���IW�Lq11%��i1��|�I�*�1�=�����<(���i��i�q��f�>N뼌�&<x�Ƀ��Gq�T.�bB�䞼_%���qJ-�!�p
U$b��Pރ�q���:�ӆs�HvϪ�3�#_�	2�`aR���ȵd�%d�yZ���5��X�C�`���3�tBC���1�̤De,�<��@O��{@.'ݣ��~,�w+z�֝����gF�a�L7Y7XըP\�O<���Н.Ҳ8�=r-��6�������*f���L!�'7�!�͇.��坚^�� �M������-��y��@p2z�����FYM��!t���_!�}.�����D�:�����V��G4����J��huD� ҟ�c,F��I���+�V�Q6o%�R��9��k�_󐨜>�#�i에�4����IH
l�!Y����U�.a~��U�\�����m3����NA��c�hv�BE�A�<��ST���/��߿�E��<T���0���&�7uݚB��i�!���N�M�(��,���뉺jh ��n�hL��lIF��8���5�I.K0�S�U w��Z�W��[rh�(_��sk��a��!=,��^"^���~{XM˽���8�NL��5�Y2�*�ż�#��di}#c�H��R�4=V�+�A2�h�/�qE�L�aŗ�@��{��
'm
�d�	fɚ�-���lnc��ϥ�T4��]ɖ�{�R����.��|�������K<�ӀP:s�%��2i���c���2	_�:_2�/��!isy���{�M8,����C�VL3_�uhZ��Ü�eu(-���<$�joYX֎K�j��KA��dah��l��`��t��z��m������D�{������|�׾�ꇃ��g����v�)�2�#L���g��WJcӋi�-�f�w0ʐ�}�+����F�f����}Wǯ72�I'^�&!u�c�#2	�kVC '[�Ͼ)��:��7L��Y�i�99a���/c�E4x�"�W�L����]d����W!�~���8����O�*~xJ�A��\ �?GR��t`í��' �tM��JU(�^d9Wg�f���(]�t��L���;鉓�P\T��m꾢�I��L����`�T�c����JEd,86&䖨�r���6a~-��~(a�pE(�p�PC,��?�z�Ǌ�Ii�S��p~	4��p�(�DU�;��S"�4�|�C������/.|����G�ѣ���{c��R/��cО��;EXUP|<\��G�lt��{���+|�~�Bզ�h�M�d�5���D$N'���~]�c�0ԯmœa�a�I�4=���'QIs�T=r� 鮴=g����U�CmVcΦ"�]�Ť���^�}7�y���."��L|�ɄEÝn|Jjr#o�>v�Ϯe*�3����=)6�!AW�Ge��W�h�sRiO$hI_zC�>�$A
�("|�u�C��(
!M�59����&9]���o�<��C$�cR�o@;þ��5?8�:6�z�8� �ƍ%"h��F�WuB���[�Ρ��01�_�̀�-g���3��w�C�8� �.��	��eN��E+�eP�N��.ܥK�3XWrkt�����;~��x��H��
>t��9��y�<�sC"o�H�������}R�b�1b��?�^-jD��-'W���N�kܻ�8Ή�M�3�88�(�R�l��J�Z�[�dx]S[�Uy����٪�Q�7#u_� cLyċI�Vjb�kQ�@UUs8��%��}k���
��A'^�aP]�ߢ����Rx�S�Ɔ�cϊ������~z�q&.Z��{���݄�uA�n��F�5�Y ��(o��b��Zۊ���3�}T�·��/�����!��jfX�DX	�!(x�W���^��w@�����n�9�_C�l-�(��Y��7$�8n�c?��#����?��xCn�j����ERlϒ�@9�K|��9%�
��6�f�s��(�#��@ovd�?��{�O@���3>w�8��S#�@�ҏ�w��g6��|��<���3L]TS��aK)R�U������F��G�����	�@�t�� "O�#N�2p��^���_�&�2:��c�Z� ��!���$s~���{ޝ�
�s��y���L:\t_%A�`�,���3y���H���%o��N��|:X)��������cBs��U&��y��h���17)�L��]w�&��H箫U���m�� .����o�Ō���h+�K�Ň�2�a ��Im�5���o^m3;j���?�^��&?����٧�1䴶;G��9�W��u?f�_܊��ŝb���N�����@1�q-8�,c������V� ։�&-)R�T*f[�YZ[O	��ϵ�Qknl�����f9���+��{FY�ш�x§�8G�>����@3���2�5jP��B4�U<G/G�&�t��G����v��"`���f��/Ʊ}���ylHI3�'��u��,��t3�Q3%_��7}��YdOYʩ7Yg���5�,&Ӯx�^jv�K�����*��x�ܐ�9�TH7 ��E���}e*d���2��RLB�G�6@i�9��������vt,�sb�Q����������)���d����?�F����:iZ���S �n5�ͮ��Œ	�Tl@���d���S�ì��ț[
&_��VLxAa���@��@��N��v2�(S��P����a�Ъ�:�3����͎"QG{c�����M�ps[^ؖ��jzLaH���f��g�Ș��_�
�LN������J�ts�i�tg����M��*��L�ӭ*�a\}2���﵅��E<�ѓ�\?��e��6"��ͭ����@	}˚;��3|��ǯMUQ n J���N��g\񹩴�ؿV=-�F[�����2\wƓ2M�c~�� ϲ�u��xר!�X<�]Wj�T�n�\��c'�?T�怦�f�߸�Y'��Q-!��Ş\��i�i3���	 |�xf��`XK٪�RS�<> Er�Bf�%{d󈝦@d�p��T���� �8s�<QO�U�?ޛ��e"������ŏ�����=��yA�8"���c7w#���j�]����gÆ����^�u��ŶS��&����n���H���wÅ9~`�X����Ϲ�R��O^:�`�ݒ��4��n�#�I����� ���g�J�r7�Dn{��E0����*�@0_�ѹ���q���%�!.Pe0 
0M�䒶āka5�X�y�Ӫ�=8�n9+�� h��Īa�C2��n,��ƍ�Is/x\��(�3��B�S�P�+��ț&�pt8�����'�O�fDe���TMDD~��\M7��+�>e�Z؉��'�Y�����7�?���`��y)hO���q;xq�M0�O+U�zS<�}4v�pLYo������T譣���qɚ�S
ʾF���T^��7��P�5Z�*����3�����pI�-���A:��,��PX�~�d�#�"�\�l�'ʔ�hg��
R���Q2������)���Ě��L�OӠ�D�Fː���ܦsb+oQoV�!�7n���o�MW�P�8Ŷ��|����eM0�r�,a���0���x��[;>�����1M0���<?����ə����x8������w8ed�P�y�t!�E'A)&��9��,�JPVƠ�<��S����9,`�Y��6���#fy?N��AO�c��5�+��PO�,�*��g�57��dO���h�0����H�ū�IUy*���x$*i�G<���J�e,W���x�w�ezz_�����:�R�3��H�ǳ��,�v5I��Р���4[����-[b�t{i��qg\��@��=ڙM�m�a�����z�����ҁZW������&��,Оx�?M�
��BjĹ��5��-J�Fe�zO�E�m��i>��u��Sޗ�Ts2�����*+��A��ZҖ�@͂��A)� wn������Q�YeSl��?7�G�醱����?��|���)�$hݴ��nh��37�L��؉�C_������O� �����f���������o�Ì�s�ղ�L_y�[�v� ���=����'B����L����"��&�eZ�
�@<��`�M�bA�T�l��=l1��{����֙{dx'��./d�J������M޷)a������8E���fUw:z���1n�Z�rW"k�Ԃ�4/�_c��B���� �	��+s�]�3��/�*l�)3�=��n�����3~D��������*AI �7#�({%a�?h��g���
K������ �6ۄ�����%M���YL-���x���G-z� j�17/�}u�(v�-]���e.V�$]W�2�/4��2��)h1�k�����̶����Ɲ���18�j�[=ʜ! + Xd�޶4�%�,����L�9"��4��&�ULf�*U�.���_�DO��1B-!�0IMa�������k웊��x��o�활P0�}Z@N��Fb�6��qe�3w֮���]/Тo� ����2]	i999�W��JʝA��F,��e��j��$|hBˋ4s��Op\���5�To�����{���4�����;�	��W>Oa��j߫c�2��f��5z&�=!hl=q�zn���`��ޝ�ۺ����r廱�������2}��������,q�����`��8-G��JxBrWt8����>�|R���wu�zo��-�e�ŀ8��zs�o�_���FC~A�-�~�;����5ŗ�%i����!��eN�+�O�ݝ�/]���Z�ɒ�F�2��szS����O�Hq�[
ו�۲���(�i�G�G��4S�M��Ŀ?��?P;3���OcZ��Z`B���X�~�hdnb@��t�o����%�#y5S~��fˁny��:��˾vww��@|T]��j�O�8>�_���R�u�\g�bֶ��S����u��|k�����~S�Ii\��PJ�

X4ܑ��]	�W��@�诶Z.�R���<`�L� �%>�u�]ҏ݃�z�e�q�O�]PT��c�JP�j��f�'�l$uЯuRebK�(�����z�G@�Ħ-��z��3i�w��� ��q���@2���bN���ٮ��'mU��~U}Ѧ|w�u�S��d��,��+�o}�t�:MQ�f������Dܙ��w�~S8���
w!�r��Ͼ�E�U�a�Wu�O����w]ʫ�Ԩڊ6谶���C�E�ׇ���6�9�!�{ A�p�_t�_(�OS��>��'C)�*�ؠ�&��_���7Bq�8p���lP�C��+���5�j��s(UP@�\��Q��&��N}�D������uy��MsQ1s�Z�\�z�(e��"X�L,��~�oa�>p+�Cv���^�#��L�u�VTT��SÁ�b!k��'�0�'�O��{@QzW��&��_o�{<���C3��bx�����uv�/�\��8�W���VD�L�`��,Ӎ�q�F�rR��iv��⪄�g��0�Ix�9|�į)ˇB%p:�ʦ�ғ��׿n9(d��y������8���ն�AP˪e�ݯ4(�iu�a���4��Up�<'���E��m�Bw��lҸ�i��tI��������vdN(��D芘��A��A�xńwn9���|�� B���5�"cp���^��P9�'O���mkǜ!TArAy=I� ���"C��Dɇ~�j)0�~6�gz1�ע�&�MiŹ(�E�u����W�(����0����K�Ԙ�"U��y0�b�^�PS�(�XZ�Ʉ���P`D��s)
�8��@���G������j ������l�L�x�-�k�⦉���yH�س��:ut�eNh��ԇ1E��n�]��2I��Ż�lp�#������Nk����ȴ��e�4���X�qԨiN��uխf�5�[�6�*S�V��*��D�yY�4E;a���#6%��%���dݥ}�WV�ƶ����-���y�d�~h~�[%�2S
r^+�:���26Ϛ#H�mV�݀v	щU�����HV������[Q�u������$"���;���y�36�4i,��ڙr1�*K����j	����B���L���V��H��P���N�&������ �m�M���G��ّU_�{�J�S�-n�޸d1ʸ���]G�]�ʾ#�	�!u{����.�pu^�&\��kTL���?�]�jmiR�$�1=:Ç������wa�E��oZZ�c�� s�9��3p����q���0*�/{:��vS�u�b�s�˔��`l�����/�F�s�+44��<!��a=+�͛�1������$>C�˗/��T�R���0���+~]֔J�{_]�k���cC��7\��a:�߃|2rz[ޔ_���h}�y��zh�z��=s1�-evI`WV(��<�����PhZP�����ƅ�d�׶�V9�ʧ�a4�{������4�%&aLȑ��#$V"~$�+��\���iX\;鷙Yi%�1[<k��6GE��F�ӿ-zęƀ��w�/?����}�X:�Q7Cpm��\�{�������޺w0:������ߙ%e�������k{a�M�]�Sg�'�/g rB�R�A��ե�%���R��7!c������<ɗ���(_�/ ��l���y�]�^���_��X���}'�q�v��+�/��UdEp������f�j�$��2����B˪�|���w�)^��E����Ө7׸��(Y s�
W��ϻ|_��,k��]*k*?&ڶ�e-�����|�zy�HO��4j��lp���ͱ{C�򜽟;F��2���;'�5��r�23���y�[�����$���ɨ�'�R�A�aC|ΐ�M��7�s%;s�Ka�\mQ��/����p[���~e=Tpm�9Ƣ�Z�j�;�~��w�U��Z�Q��N��	��`��1��/��6�5����v�	z������~��b��^��� Dr~ps��V�뎆��R�mt���޷+A��Qs�n���L8����(+���VsݺIm�|��c�͎��W.�L���-P	�z�5W���4ۼ=f�I)��`1�8�G���إX���xJF-LAp�Cř�O�ҹ�,���w��Ս�3I�jy�jy5j-��
�z�4>_н�!�T�0�7�t�m�b8e��ґM��ԙO��:�?\)�74�/jx��Ӿ?#y��ӳ���&<�����+q��w�=_�4��Bʋ�H[�v�5�/��:]ԑ�G�\;�{h��p5(_#	r�|RE�i��tW���]:m C;s�i4�����_}�Y]|���$��bL"�XʉH��&�oC������yW'�xȣ�,��i~�c�*�I<b5蝬�	2�!��uut���w�jjj��M䔬 �w�^���U �Zߦ��+'��וxdl9�sF�R�	_�:q�郪95W&�ɓ��.[��0���]{x�!yx��),eݟ�k��N
�����3-�[��!4Ut�Z�R����d���_⟦�D�����V�~�������A����%KJ������/J�T3��Y�Qy/��OxR{��$��1��6i�r�U��6T�Weg������N���gh���
��`]�[c?���1��rCf�[�+4�����
<�g�k�l�V�5G��8�l���{qwm)$+��xk�N��$�b������ �����Ԫ#M�x\�`@,%�Z�p�\�n���U�_ާj%"�<��}���~4q�7VvK�N�K�xd�§�KU��� �)v�G.��Kբ�k"����<�xm��j0��n�� �F���@O�<�5�:���X���9���ꝏt�Q%�f�ϫM�����Ցj����O�m
*�L
N�B�Vkʃ�?y�(�r��δ��tJ�\�cAT��� �h �^�Q�$ꙩ�^������Tt�C,����B��e��:���ꐴ��[�G��Ȕ~�q5���U��Z��P�w�|B�f{[�$��2�+��n��O���hwNs�r���ƣ�Uj��sgg�I;��-�Qh	H��}�eh(�:\=���ϓ��*�
��s�, .@ޢ�G���oO��k������){��c>�
��w̭ƙx������P<,���1��<nO������8��a�Ij16~���_��y�/�$:3If\?���/�>�<��u�B�ݣ_�LR��� >M���6}�R��݁O[&�ꈐ�!�=M����|M��}���v��̕<m�=�/SnGV����/���/<�9��;��;�+�s�����*�s�s��c�o��ر?�� ��a'��� 1��c-I+���$5�k�/%4���EMM�P���:έCP���4�魵Q��D��l�˅"5~4\ވ��H��GR�&ISh����qt��l�o��(1Z�VP�UDզ��ݪQ���Ԟ%E��������*EEQ�hĎ���{������<�������C�:�PaRQ
;Ձ�+\ ���`˴��-ӄLL���@v�C�C��_�YBR����g�g�\7��x߂����Rՠ
*��$�����~^D�fW��S�w��q�ܺ-�Hl�_��՜.k�%�A�К���J��~ł�$+kl����b^�,���j���3�A' �=�z��}
�<�����`)G@��3|U~l��(3	��|1����y(�g??y��r��roº�$+X�J닊��Vn �`� �6~�5����k�B��E�&��fN�vyFp�U���`,(����<a7�-�9�����0Gʸ���|�#f�L�2�h`M����k�(~��@G�6�V�d�D��1埢c���m���!�0[AfT�BoT��'܀��"�+�xd7$*���	y[�2D-;C�/
��I����&B{~1(Ӣw���~KF�)>�XX�{�F��k��i9�|4ӀܭfMK�y����!����X:MJZ�xVE{�.0P�o'�-%%��X�u��[�"Ǜg����-�R$dXj�1Y�tml6���7��0̠�m��h59�._%W�9�⧛[S=���#���v���|#0t�,m.��bɺN��lX={��e�x7�2�t
[��|���|�C`�Lߎ� ��������B�N�".�%�� e��<,���.��/!>ڕ�`U}�##�-��_���O�Zv5�^/tC�aY��4��l��ã�]����ˬ+�F�:�j`h�2��x�3�v1�w�{k�k�/l{�9 �u��r�>�c���>�ʻ���S�J���ɹ�:̧�O����_,���l..�zq�a�S����5��9�`�ج�]U*�o���=Hv�k��2���W-�;NC��B}4.O�91�)I��JԵ�$���3��R8.z6u����2돢F����?� Y��2;�͉@�"Ud���W��?���x���hh��� ��:�Z�|�x#aur�s�#)Y_ήz��t���Y��v����U��$r��V���� ��?�Z��;i�J�	����줩K�I~/cG��q�r��rǑPH<�宜D��߇]������REk�w�)��Q����"�*���ۃ�=�)"�70� g�cy8�Z�I���cn��*���P!�����y�8�7<p�{�[
(y����Xi��ǈ�&��s�O���m�2����>�"��0OHbh	�%q���b���=��������)��ؘK3��m+���:�M
��b,���C͘v,�L����
��O�U��%̛��Icɾu�Ɯ���P�P�"d2� n�:(Oi�pF�9{��9��}�
����掼�.
�~��o^~�C�����=m�y���0P�[;��N*x��M��w}��,Sw��FE���P/4��,s'd��m���s{?0~3�b�V�z�C6�z��	:Z������q�Y��gY��S��w?XiY]�2�=t���f4�׮�J� ��g��=!&	dH�ގ��FJ
����D��7�OE�!`9x/���X�M��v���h������vW�i�ьM�.�"���y���R)e�����=��˔�H�W)�����R����m���H��4���>(�%>�ub=�ĕel�kDc]\c���� e��|<�uB���a�o= K �5p�S'6\UUӈ��1�7+����I�6��>٫vz�nh�T��ה� ���b��M��8�`	��th��`fb������q���;�b^���
ĭl:�(�+�,���ѥ,�c�`/�P��b��r�Σ�����5��܊Oxa�Oiw��F��� ���P&TO��16�`�+��U���ߵيz�׵x��QȬ��~�A�^C�f�"Z��3��r˧��%��cXmqV��q�A�M�rE�m�b^��U�倭�0�4�f�]�x�r(MC�ؓ�/h�-��'`�O��&6�/ǫ���N��,�笻��mTZ�f �NH*֦]�6�*�b[3��8�)ƚކ�q%�5V�O��g�IQ�Q,�c���`_�&�n��r��� x-}	!n���ezVo�T�SL�*��Ev��v��b5�^��Q�YI�$U䕯���=]�:��:܍M����Zld��m�jh��=joqW���h�I��G1����y�~��c�ܢ괍��cXǉ]>R\,�$&&���F�v���z���dcc؎�0�+׭Pk1�<.瑯l��2녴 ��f�'gD�
����i�/>�d�QE����l��^Y�����,���8'�nh�D���	ϩp�mr��A�("�k@o�xIU�`���}���Z�Y�
��:�`��j �ÑtV��0�V�yn����	⢾�_E��� Ԫ���/P�͞�ɪ}[ʶCn?�6��W�f���q�P!�v+=;*\f�Gފ�u�K�#y0Usa�6�����	��r)�Ȕ9"ؔ���"�-�>�����&��p�8*0+�;���d0Z�wP�%1� �'�F��J���Ϋ���1X���!~��{u�m�ʛ�o����t6��C@��:m펍�$�0�	 X�.�ؤ+IO����u��,c�/&X���R�@�Y�?^S��K�!ހ��O|-�|,�K��7�K=��96�8VO*���<�߰L��cQ�d��{�o����Ϋ˴p��ǻ�g ���΄L� '=�xIO#Idy�M&Ix���z�fJC8X<b4�s�3�QW��]'M7?��RK��1�T�p�G�$Vѝ�8 ���B|�o���2��y8���k�1,���09�t���`����ǯ��Ì&ħ����V��۲�o�#��Y����	��$}��Pg��1U��i���J��̫i!����N�����L�e��� ��*Az	�l)�A�.~��i^¤���{�g��#�?.=��`}�ol�p�y}'��� v}[[��:S9.�}�ݯ+���wo�����/夘e�UU�[2�y'5$���D��;Y��q��|_�6���`y7����XWH�#a���xw��A�&_qx����Ŏ"_�n�hg�c�>�� f�͚ �$�٧�/{o՜����$�\d F`�z���
�����_BT}][������7���t�&�-x�\�ì�v��	O&g=�>����V;?�0 ���{WW�R�� ���WPիq���^�-)�;��D	���i�։���bE.�³ 
^E���#޲�zk��,��\�L�B\�q!�\�2n�(~�\v��L�nTO�9�{6�UҌb%y ���O�N�K�+O)�()%��l{q<��r�􏜔Gw㹏�~�9Y6*��������E��}]n�)e�G���INaq�o�Da����֍	�t�m��l�o�)���U��.���[�A�];���Y�"�(!;\3سAP}� �.ԧ���	���цK�F����.���:��������׍D�e�Y1�l�z��P)�`�l�J/�����k��x ?�Ij�ho��5�Bqw�_rU`�Z�f�f�N�[H�3��>M�5�
�bkٺ���T���f�l�|߿ �_�o�`�����PW�������3�%ʀ^d�N"��ua���I��'�-�s�]����A8�+ʡS��ҪK��UQ��1�g�����2�;Eǥ���_"*\���5����p�,�
1���r��o�ޟ=�=t���>'�w ^�RiX���� r��-���Q*Bg2T)�r��r."l��:bw��vyL�k�3�-����D���=���� ca�!��}o[��� ���P�ϲj���"��00���`��y�l�m�ۮi����4ֳ�ORYNA�Q?<~���y��0+�}�y�脮l�o"%��%@�d��6�Z��+p��"�V9��6�ϦD	 �)�2Q�*�^k�Ɠ-��?eP8�i�ˆ7c�2�,YԀ{��Y�����C�@s���{��8o� ���{����T�V�b�!����݅�xN˛�M�/q*��-m�it����ں���B�l���;�<v��թ��$��߾9�N�0���8?6���~Dރ۱R��o�`�����y=�����>�V�zL	Rn5Xe��tNA�0�I�8I��l^�c��Z��Ʃc3r���_c@�,��$pT�����$���I���=N�`]�L��m��"�jO��D�n���G3�%�~w������l�p�J�'d��!�kl\^�ɧ�ְv�\ok?��JW]5��T�u_�?{��8p�[`��N:]kVz����`Cƣ�EŎ��pz??�`�:O
�g��s��z5خ�S��߳�����I�<�*m���a��Yl`�;�KL� rԈ�]x\j8ל��n,Q���Eb���h��7�"�3�Qn٬p�4!�)�=����y���v/u�ux��aJ�W��p�i��W���֯0�m����%�(�{�4ֈ�HAVV�χ�,&66��?eQJ��211���6u�/Γ,���i|I�KK�:j=r��Kl~a"�H���	���e�7M����S�ɩ���_/w�g2d?!q�c������o�\�V݁�$8�0@xOȨ[I��/�df=Z�s]w"��@���*jg��i1�)�	,�D����u=�1�˃�Bu?_�t�Ջb��H��Sm�F��
�)�:,��-���?E/�:5Z�����lq�՛x�IeX���R.X.��+K�TG	=�:+�I�G��U�h��ܗ�u�����'��#׋��	�[��r�a�MSq,R�_ͫ�E��L�>'���+ )B�!��@�v���k7���2XRa�b:TH9�oz�����u��߯F�"��2!mf��ԟ.c��A�0�n�]r ���3+�+]�e�W���q��o/f��������ΰ�(��R`\���m�=M�ݛ4�nvo���hW��G��t�Z�3x����jȓ�
1���%�"l��C�$�~煩�SM��ϙ���Z�9���ܼ��||�.�V���ў���q�����B����<���f[��I��H�.�?�]^ԅ�1��N�;���)�n{�Y*�PN��)@/IOx���v�8j,�=��`M2�/���^j�]1F�ć�g�����A7��:���5wʻ��q�%�8����!�%�4*V۲���Gc�Z���6N'��{Z�UQ$��'��۰���O�ao�r��Y�"bf6��m̀�=��Ke#��y���Q���0�%E�r7��`���ao�[1͞;e2`MWz��r�����j�"��1j����*��?�+�.�}��w��`b���ۍ�Ơ˿�S��x��n�n4� 6��566ˡ/�텳;�ݥ��&���K�WgЇ{%�t�w9׹�{�e�1,N��QPo!���DDº�&7X���mW�d|'��_TJ�<�2�9T?��e�N̖�E��u��(6:.��6��t�ڭB0x�֭���&�0�h�ca�Ln'WZ,l�c�UC���*+����(i�^?:9�~*�@|�!&�����L���*��d��: J �}������������/�ʳ������D�:���!#�%�ꩪ���YYE6Nn u�/{J��V�Xo����.����o��F��-�:��6ˌ�7�Ƌ������`�2��f��8(.��P6�n^eH�T��Bo�Ǌ���TO����X��r:\�uAO����6���j������'���鼺<#�^���{Ls�7�0�zں�b��M&lvN^Y���XQ$P���/r�K0|E����ⶄ�_��}���� t��K��MؠLk�����U&˻e�\��>�Q��姻�} 㪧���w�r����8�="g$]8Z'.>B�d�{�'��
�O�EM�E}�X���p89�;��yr8K"?!�Ab��ǫ!��h�찪)c�g�\�JY>펞��2"A�=*�X�t2!K+SX�t��q�^���"s�D��ڟZtS��d%l���_΀�(a�#�����le@^
N�M$wa�8�&��@�9{�P���|�٢^-=O�`����PB���_,u��W+�'~�bܞ��U0�T���ɷj�8yz��TN{���[�7F�k�T�M/sc�
ߓ��ʢ �h��:Q��j�_8���TD�[IY��x2��Q���}d�b�/����,�Ì�V��Y�K_D�; E�de��\��앑6�r�yb�~����9-��n6�C�v�$���/44��om-����qE�/(����n-��}k�1��GG������vv��-�>�V��r���DN����?CU��K�ѥ�FC�k�7��Vp��(�T�&�M�ņ���߀�Av�ɏ�'I� n�e��l�6�QDЉ�]8������Of�����;=�w	��Op܂���:��G``e���r��"�U�cƭ��Hwg'?�O��:���s�Յ�7�\Rv�o�t�+�Р�#�BI�5^�������HՀ�Á��42�9|�j���Z�����s$M�������1g60����7���I�C����,����\٢��ul���I�����8`�	m�X�fMDG7p�aq�-.��E^��!DN~m��vۘq�`ž������հ"����қ j��vU��H_6��~�3r��� �]|�<��2{ez���K2��NB�m(���^�s#!w��:Lt�U�u,��S�d��T�5Έ��c�K7�)�U�^��^�5�Q��|z�`�iZ��8{?��NyA�ų;Mt*+f���;xP+�W�y�
T��~���o�Ba���mq ������ļ�'x�`.Ч�}ww�/:�	D��ױ�C.���%�/}'��2a;�[�j�[�ut64S�e����<��^ ����!���)�Ͱ2��˟�c���)���]��<{.n\$�'��dZ���Y�����QX�C��v���^E>�N_�ئ-P���}ϋ��� (E	���_����j�&.vo<�
��M��ϛ��DT���5�XZ�64���2�I��͖��/���:|w�ca�6�	�%���M��|W/��&��~\��E�D��b�+M�U3$�R���W	��w�x�z���g/v v�#��V�'���s\v�E���ft_��"||r>r�W�R7�>"V�4 7��^9�F�TG33v�T�ꉉF�Ҿv�jq�S(��dF��x��>�յ��Ҩ�����,���[�������<[�j��t��5}*KrZ�:^p�۫����x\�W�</�����-�<ʻN��[�'A�K s*	-.Ew�5����3��p����K�V�Mq��Jk���M�8?X��|��U�ZЈ�_T��yōłlm�	i��h4P�NÕ]00P����5 砑�4��<�~iP�����@ʻ��W��_�=�4A��<�jW��^:_;x�����-���3��H�%^��zI���%�ug����ƈ��#��=:����-˨0�oր+��a�-_s��m�:X�OM�ӘMCN�M�6�~����ټDL��w�~������������D�G3E�!��\YƐ��*�
����kk���w��� j�?_8��xi���9e؛������Q)����H�V����w�nԨ�Y���J�m�k���}�i��͋� g[��Fق|��%[��7�ْ���-��ՃU���:�����@%mVو3Y|n�Ǆ������5q�����6C�^�q�Xi]`��"������i˩@�ƨ�)	{�ʉQ�åR�jCQQ�����
!�m�(��[�Sn09`o�7'���S,�Ύ��G��.:t��F����; �mn���Q/��qh`g>�����]�o;^Y��<��Wؚi�֏[ԉ��2��9L���ٰ�jn<��-����t�\t��@j�mOd�.���!Nw��w,���t'@ܿs�8�.��3����8KD�!�/fv�y%:`�NV�3��r�1������V����!h�ġ�Թ��b}�S�����p��uvk���B�(pz_�^��]�8��$qju]%���ˏrpj��W�to��]�9~-�qܣ�۟���޴��o{J��(Ӆ]���k��߉���Q�Iϝ5���@zd����)8Z���jg[�<I���6ͽ~4ﲅ���}�Q��@ћ�Q��C�����M|���ܞ-��kL9�vy��S#�EンF���%+�!�L�0}�:t��\����M�4�D���_U^�������\LB���C�(PT=F� ~h�|OD��[�a����?�(�e��Fxb\i�>9(M����Q�{u��jt��	�~8C6��j�Q������ń�-�vq�E��S���o-�:1ֻ܄y��W�҄��vv;��0���-s�J���fsJ-������pBuuuB��G��#��{�S�H �z�|�����U��^6�i\�b
�x�L.��5m��w�#M@���(!ݧ�|(�m$}`���6��	�\
��"l0�bs���76���YQ�`��6J+*�`ƿ��ǉ�oL��znx$6�^�G��U�H�G�줭ٻ⠢xՅ������P��4 ,:�{*�/)0ӑU�.
:�jq`v�7������F�Q����us�D�7�\j��grBk���BKBZ��Q&���;���'E�4�%C=�GycBZ�F �T�3Ƭ��_��征Bv��eJ�hB�}���;��
H��`]6}uL�Z�:�"�pdYHqʍ:�݀QQ����n|4���Ԃyx���T8J�,I:����^��y����:^Vehg��0��q�L��AI4�k�W�F���4���uY��!������-G6;n�R0^Q�~��a#�}�zHT#,ř��h��2|�A"��,���Wԭ6����#7����l ���b��<��7��d&�c��␕��=���`g��9�"�h�nY�pX�^N����ֶ }$"/  cbv��Mh����$:��FF1ۤË/�ˏR�!ޓ�&��1Lԉ���A�W˝�Z��-���m�7LkC8|xcH�?�
FWB����qP��85Jw�oC�X:Tb��-[���q�����32H���h!Hu7�����|�o�� b4�u]��c�%�O�ͯ��uf��|���{���o�.�䆟�kL2B���ȶ`��6��?���䣨G�����/v�d�����2n���6n����g���� �,�w��e�x�I��<!lmcC}qLK�����?=� o�3��q7��F#wDX��է~G����2s������nʻ��H���^���{^݅0�!WK��oԪͳi�z7U��Q,h�o�Q�)_�G:7�P��� ~��$12�W�W�D��:
�����A�t�M�
_]|z�2����v�l����d��fk)�'���_gi*�(�~��V��W����ߥ��A����7OPP��8H��U�J�,5�8�+��]:�Q&�7y�xv�E#x3`��#r�@����ϰ���g�JYm�en�-�ٖ�4���3�K�H�W�u���IzI=g��=�9���nwN�U�H��&����:�h�Iw��.��G>�����c������Y0�p.c̴iEM�Tg���T��Dt���)�CN99�#�I*�=F��E�c��zS����hfRq����S	�/=�jE�KQ��F�)���Ob��l����Z�M!L�O_uɢ�,g���lʚ�NO�v���6AV��X����������C�!�B��aA~)�\�{�P���\�ƌ8�{ҶުV�N`�'f�T�u��������#���Ȱm�[����h}�A�(�R�E�S8f�h���Vڄ?�Ke�5"[�49�p��Pq�a���4�]u��}��J�&���dtGZ^�â�g�`0g��½/֯_��ӡ�����aH)��;�E�5R5���q��:!|����.���-\�<��Yx�����}��9k+Ku��_԰J���(mr�Y��l�^'�뵢��9/���9�� �7�C�h�.�9&Z���[,$Ѡ4_���i!vQ���'(��� ��{�c���	UIjb}�=W�ҳ��:&&�ti����(�5)�9��F�8r���Z����k�fԑf�Y��t4���/��lP�O�?�M]�} �}���+E�z��U�9`������$o��`�оT�\�<���*6߄mFi�<|z7f�+y# Og�Ǟ�r����	E�����}1'	P��f� L~Ym�'�KM;����pco��n�!6����p_!���p�@Ο�p��r�&�)�}�;���ѕ�N��V;��Om&C~�m^umt�(���WkK�T̃ju,x���Ϫ�`$��A`>�'teH��4�6�Y`��k�K/����kJ�ů%b�hA�%��r�m�c����S��vjL���'ܤ>r+P��f4s7U�~&��c�����Sy?�u!vb_$�K�l֛Xa:O5 y%6KOW�}hԎ�'7�%���oN�M��4JY`����]=�mr�eI����W�����r�Y7.F��U�;ʗ���(�({�*b���Q����,i4���)�8��b����F���T��Ü��]wXx]c�;�xe��Fq���Ix�g1{>�#����y�ɸ��ar�O�8�,Ƒ�9�)���֝ZI�?�ܢ�2�?�@,���kA	kQ�p�%�(��y
�GBƀ���- E�v�0/,��Y�^��C^�3�x��V9n�ha�nGv敒:`�o�Ud�7b�ы�����@}P�`%PVv$B-�Z\Fi�� �njb-	$>�ˑP��F^�`�}�[�X�2ǹ�aF�V�~�,�>�,��*5������ڜ�= � ��o E;�8�R�V�{���s|��JޡF��7y:pۚ���sV����k�Z���7����bm��ĭI�W_�G��h_l��`�)"�W�+�Z� &�I��%����y�,-�[���f}�,�(��
y�5҈�*��%}��qL'�)�D�jc��ץ�x�hw��ʃ�����&� �D�{6�������?��:���mj��(��6������1�� �+��4J3Y�d����[!�&��A�ݱ�֜"���F���2veA������L�Lh����9�����]C���v���0��[���,$�!��m�T ��i,�!���#<]�q��_Z𶈨ma ʌ�xz��0��2���4�յK�����ۏdyd$�!��0xrC�]���Kd�9Ĺ9�'4����s�y�����W�y��&@a'b��#"��<��46>to��T`(��\���8�q��ӛh�0ۆ�)u9Cbo�K�݂/.!��߸ǧ �S	g�=�=ƍ>`�����QWȆ���>�Y�(���W0�3�\0�ai�}����c���f�
jӨ��&]�w���p2r�	i��1�ׯ_?z)�h(�%dc�/r��sS�C��(rx�W������c<NQ�"���:������B�-�������;�*Z��x<�p굿nE�~L�Cg�����`t��7�C��`���Y�7��Ǖ��-8ٔ �k�[�/D ��*�#n�����_����+�fg��|��p�:��B@�@l�ް'���/c�k]嗡^���:�ƅ���,���'��ߤ���~w��L�|y�$�w�(�Q�|��P0��J�)���2v�S�f�݉2�1�[T��F�����ab>��J6\<��]3	��	����!�6܀z�����\G��ϸ�5{V�-�h�*�˼��A����d)V�w�����5�6O�E�����x;��(/�UYy팦��2m����od�G�ɶ�D�n����|��|��#;�Q-��5z~��-9��͉G�ɼ�#��Y>O�g8������h>��N҆�1�n�=�����TH���2)h��;�/Ŕs�J�e�4!I��M���}��텋�m���:��x�x��k�>��tHq�F՞��Ѐƀ�yd�w���-����YLF7!�aur�<#�}���>�ʭ.Zu�9,N@��7ģ	��I�\� �=t��j���TU�X c�00x+���<�^��@^!	 Q�1��%��X���;���.>q��t��;����7r�U��MJ3X��n���Ѝ<�WƤ5N�P	�"�iө�"|^���-���q�Ẻ�v�V��'=*�_���4Jr�N=?P�@m���%�t(R,3�D�����7c�Eᚐw�r���Q�,y�,`-{�k�bx�=4����Yw����)����~aP\�X#6R��kđ(�0ґLZ�"Η�\��\�|g�s{$'P�����k�p+UQ�<��籃o�	�%��,:�<
��uv�R
[3�2'.�A5f[��d	�Ի:���A#fS�b��^�m�����WӬn(�y�;�.���u��jW��K3 ��r{x<dA����ѽ?��?�k>��er����i���AL3�;`g�N߉�/0{�U��Vζ%��%�W�/Q�԰yΣQ�D��bS��e��R�l`���|�[�F3Lf@n���<��G�� ؼyα��G补��HR����wD0�B-pj����V��V}�3a~v�w�{�%r�* O�+�-GX+ͭ��g�����#l珩�9C/��?T|2<EE��םۺ'|�O��m2dw��N�3J����[���g��,<L;�50��ł��Xa�V@	 H�G��\��a�1ӗ��>�]�ac��0�U�hC1���s��J5�#�]u���A��p�F�f-�"o#�|p����b���A�e�>�Ֆ>�Pn�����K.�!��(�E�� �����$�z*N���;[��$)�B5ĩ�*lDo��)�ikh)P\p�����H۶뫧�[m�X��a����:	W�j�㾎����i�Q9X ;�!la���I�؍�n||�؅K9��{h��s"R��cuy�� ��e������yB��D�%� 4��p%zN���?fyF���=6ǽ}�D�Ʈ,��x����;��)o���y�)�٬8A�Km�,���e�q�}m1���=y�s06��ϐS����fk���u(�o��>���Tv�G�~@s:��3�k7� a7��S�]^�&�q��	�J�2�&u֤c�0�b�W+)F���A�B�x��}q���rrɒ��l%�iK�9��"+�m�!�W�b�뽢�N�0@��������q���ǳ�/��fѹʁrB~!ʛ�FhI��GB�>fN1����!au$�No%�R��' ����:�A�׆�%���N�1���r|�}yRxu��!ђ;C�L珑�6�q�9G~���W�6H7FP)ޟ/����r��g��/���F�r��Ub�� j.�]��O�� r��4�[ن���ޕQ;�	�/#ܐ��������A��� C=�o���n���m�E-�i����[�Xcl�g'��]�O�d�{���̘:�&�^�gQ�  3�c�XR�1�"��G�[��Bm�/䒘?�f �����|�|:�ݦ\	J�n���y�ӅX`�;�`��bC�O�ae�p#D4s�����K�$���+�����k�����e���E����h��H���4M�� 6hJ{o������Z"�i��̻�ޞ�zq}57j�*ϛ���T�d�d����R���5��nE$ ,�������E�z����AU�i���l��^��y�]�V�ǘ�}��N\
΢#�F�]$�BR�-�����MF~�&v8���at;���,SąUMIQ1*Z.��J�E�l�]NA/"��TBk��A��~sC��o߉Ce\�����Q(�����[G8}���?x�����vZ<�ǿ�����?��r��)2*�)�ʃf�E�~
�>^YY988?��p�Sz��d�2
xz��n�0"y�[ZR�z�*�ƞ]&��]���f,֏G���b�8��M,��\��b�T���rO�3��i����m:����F�z��8�4y4Z	�`�~Ɇ�o������ޑ}1�	]�"F�ql#)O:���>hB$�%�e �Y@i�R��s�[H)2��Q��l,��˰`��HF*��n�CN[�L�X�����`*�:��|�,�E�;CJ�uvS>t<I]�2�>c_`�qݞ��VӨ�l���G���n;҅"&_�_����'�!i*s(��XYZ�����!��U�iB*���kj���{�_�N��\�}ɻ����X�%ÓL��?˅;��f4�.T�8H_�)����҄�4)�:��Y̙������.+��y���e�k�����!1ˈ�BOH*��bAн���p̸J��f�(�Q�&�E�jl��ξi�꣱]�_�SdcF�%K{�S!ɸ5��8�I�U��!c���GFF�M�`����Hs2�G@�G����M3mz�*��ɪ�Q=����v`��"�^�P
-��>!�;����>�̒* �^A~�lQ~�HOx�G�����b�y�h ��O����u��[4u�1����33�mt�i�;h9E��;7�C�>����b��Qw3�G�ݹ٩����[ ��K�O�u5�[����?~>��ظ~v��Ǫ35!D�%[B��	)���1�f[����A+<r<D#��qyR� �t^s���k�C
�� o�N>]ZZ�E�_-#���{�������G��j�z��+u����/f�z����k�vk4��ɦ2�!ꏎdVԀy7]9�1!�$s�GC�S�V���ؘ�!;:{˟�b�݅�R$�ˎ̺���'�LJ���cl�;�H�k>��&s�1,bSb��%`�Q�vy�֝N$2�M-S�ע��|�9�ԦPz�m\ʵ'���#^{{g���q4$��4.=9c��d
�ר���}�M����*���{
��d)�g����q�Y�=�j�^�L,Kw�wZ͠�!����Ӆt���a���;�n��{qG�1�l���R���S,>�����m�̼d�}���oK���+���m���\8BJaq5�C������>�1�fAN�Q�Ư�`������Y��Q��ϳ.�t� ���u_W��+���p�s}�~`��ՃЏ)��g�d_���D}������ؒ��i%�菪�ܕ���P���*p|��z;��s|6�##��&10���5Cm��±M����~Z�}VR��B��Ն����ұ����jWI�J�6fd��	�p�P�>@P��9ɗW����;�*vyY8��P�E1tE|X��z�QO<��z�w��{�;,�5P��^�v�+�<�)�:�~V.�z����]���e���P�!����k� �g�>)��>�=PI8�V��qz��������\����l��;==M��o�du�5��Mf�T�	A�8��_�����J7�rson����N�?�XF �/6��2��hL/-��jQ��n�{3��ޮ�(��a��|���1�H|3E~��5��\	��ܸ�	�M���R\�7-Nq�D�����r@"����T�����2��8C����}%�6����D�o[�WGQ�M�5J��v�2�ݻ��3�w��i�G�,���[�'��(��hTuCC�>����ª1'�������N�;���oO��M(1��Gn �p#/��,�Xܑ*G�&�p��H�P�ʽ�M �Cݎ��RO �d��9��S���u��>yBW3�(S��N�"�ah�3v��%s����,y����_��ݞ�r�lIj�Ah��y᪨�����x5�1�]&�6���"��3��ܴۛzt��36�/(�ѳ��ܞ���[��):=ϠEg��pȏ�+lK���[;�d���g?� ���T�v̙#G1z���p`������ߩ�)3�)�����k�A�,��Z��x񄶐�thv�F�-BwB<�	^�n|z��k�dnAYY>�������|a�Q�KE�COV����&gzQ�r��a.�[��͝��ck��r!�O�MQ�ѱn��,zU��; ��[}h|��;6Ƃ>��t��"�J�l��� W�r�B�N�i<���}�E������Գu�:aؤ��[�����*�����[ 1Ѻ� �bpܵVS~ސ��8����F�c����u�AM=�EE��b���ޑБ^��!��{B�Dj �B("M@��5_�4������sg3��?y�d��>��9g�]��?vY��y��WOX���g������������eɭQ��z*�5���=�OU�����6HMC����Bk �r;^�?�`�m�x_6|M�Ԛ���ꙙ����'�%����o�����Nc;�?�qL���L�|��#3�-H[w&��r~�CAg���9���yY/ ��#H�J�5�9�A00���2s�H�����e �ԍ�b����
��Dq�|�\è)yܙ ���:�~���nk�5{�j���7�i��T]��`�@�@ޢvTg�*��^`6�(�ə?�9�NE��%~z*#�z�ean��l�t.,�q �1�NϪ��Ѣ~�e� #�ӹ�)�x����$ru�b�z1�4�ld_�\Eŵ��V�럻��-��#�$9u�48��S-7_	"�;uz����'gni��|t�b�3{�X']N��'��߿�N9(_-�].fv���x�+�ދ���x����y��f�L�x���`��
��8��,
Ci@�����PN��bR�/� �cY_�eǟQ���?c�ʳ��ӹb@��*�ZOЂ·%H�64A����yZ�`�/�����n�f���2`�"qfV�TG�������a0�L>bw�4�ce����W���+Wh�Ãz&c�r���:�~�0A�d)/��Y��F��z4{���β�,�m�3d�M��{�C^/�x�����P<D�8�ث�®��j���De�A�j�w�wu�Ҟî}��W�W&�gӕLÖ*���������@�γ�P�T-��v����X͌Q�{4D����`�������crKJJ
{bn��w�χ�%�t==2�/N|����S�#aծ]��?�&����-�2L��nLދ�Y�:�V���`�<Ƕ-�3�j�w��{ꈇ�h_z�4%�=���
�7+U�Y���#�}ͫw�V�����SM��}����K���1r1x��I���V��ՠ��dm�WG܀��) _��dq��@+��N�i�S�,.ڵ�V�������^U�r"$���6}ͫ$�w�<wh�vp>=��>"8�K�������6MM���v(/3#�(o'�6/��=�i߫�R'�YJ���9FQ����X#ʶ�<x����0S=DB&����3�%)3!Ϡ����f%�]�����0Ǫ�m���}&���."�SnR�,�
?�mπb �`m#��>�Y[p�f�\!5�o����4�-:qb�ߨ^3.�f�"]o��H�R������1�=gyu�p�%*�}1��)w�R�����rv}��W�[zU�x�tk$<,,�ҧ�w����$F5h1��.>�G�P(6Ti>�#v�x� ]�Q������V0d��L�b6��#�a9叅h�!�Z_�����h�v�r�^�m9��5���<�?�<���&H����$ۺ(p.�{1&�$�����8\�|ꎏ�8Us�w���N�c�F�ޗ�|�g�=+�)����gj�poPZ*��[��ꉽ�-���1A�q|������y�u��(�Nl�Yd�'���wG+�g5�����i��e��0�6��� ��ul���ݞ���%S��6rA������t;S���R��q8j�ϣ����.�(8Ь�mP��͌���{!�x�g��U`��#�-vt�k��p��R�?�7��^l���\�{^yս<^��vGM�����
�]���Eف���%Uc�f�b2y	b򲲪���~^��Bh�rix-�eK����p�'8hZ�H= =�|(,�jDl_#Ez�r'�W/������J�������{��Ɲ%`Y�_\@k�.O�R�����XXX��2��5�Y�k T,�CK Ry�1�쫇�5`yzT��1�Qث���x��\���k2���)��l �����E���/M8�n����+�����A������Rb넛��}/y�K��O؃�8�-Z��#�|�OƢF2�����3&4\��*�R�b�����s���	SXA�偯��9��M�!�/���ؓ��������~1�8�^h�J����$�ζ���s�U�2����%E��! 4���,Y��]���z�n2�z���#��>��.���9�u���Rgn�x5h_��l[i�	�O\g6�9m_�ln���C s����?�0��s�S�^�n%���nIh�?O�NP����tpi��xuc����b����C�"ia�f�7)���-�%��,_�U�9	LH^J
}�_�x�*ub㩫%7ⳍ?��^jaoo�c3|{�D`иoѦT���F��e��X�J�L;��Ή�?}�HZDI�k%YS��~�0��X��ţ���D��pq�x��NAppw��?L��LK�9��2.4��y�'�¶mp�:_��2C��������<�_�,�&y��E3j\����ق0͜> Cv��h11��
���>68�w١ݒwVC�A^F���O�^1�q?�<����;X0(i�q3�n�0J!�j� �p�5�
�)Jٓ����4�w�7Ӆ:���-ԅy f+�r�8I8*�H�]����V��@Y�K=�b������dԟ��mA[m$O 
��d�b�)�����y��X������Q� �&�������	a��H�(�q��j���wK��~�T�1wyw��&.��%*�_A|�E\������/����xu1'�?hFc�������v�܁~@�0#!#b�ϩ���Й�3:��W�W{��Z�ښ4�_X ?93	*�cՠw��/9�lt�h,� ����4&ߐ�����O�����t�M���<j�Y��9䃤�u_TV7,��`����Hl�sN)蚃sJG'TxL��r���9�~��&N����,��wJ碄~v5sb�B]�x�듩2H+(��U���[M2�&���ҁ���n������DM���G(o0X��gKϘ#d]=+���:��}��o�<Л����ı��1�d��s�)�f��K���<Ƣ�(�Oچ����i���@K/)YiY6=��5;4W���oxp�쭵�I��da�,���--aS������e���bC���k��J^cV�6όl"%�\+�t��d���*���
�)���c�v����j�,��4}�'@�
������iX�䇿��Yj���L�
�<c�8�YuFXd,��e0�xE��߳u�O�W]�Q�eW�
g��sN�^]�K���.Q�+m���n @H;��K�SK��P2#� o�o$k�2��oa,�n-�5g�vW.��8����pl�~�R,T<�� G|�$��Oz@;�W��|>���{�8h�x������y1�w!���z�����~2��>�c')�3�M�I���O�bD�M ؊*v���Ҋ
2�)(����Ou�6���!��9�PH�)�@A��s�W)��#7NH��ʘ��*>��}#���$�N���p����D�X�!<������Ϋ��z8����p���י^�)C��	������UT��̟�+�Y��*��08C1�X����йˌ^���n�m��ύ�iC��J�����;�x�4Ö�g�RE�!�-C�Y����F�z��ӿ>j=��M���"���g��&���MGn�>:Y)���̰��~42��F�k��[��i��P��k}�D�}O3�+���	+��<&�ǎ�k���&}-�X�B9����x;C��l��\88�A��W�m���П��?8`�b9��TZ�~��-��ee�O3!���jx,?#^�ITȋJ9�i�!�>z	ri2.���&霣�c������q�Q�4ט	oGM�a�}SH9u�Щ�"^�J��?yaeЍj��%�s��~&��j�s ۲~	_/��b�o�Ԏ�8^���M+���䝐�\�L����T���4r�Geq'Ar���JJ��}ed&���荓���#�ǫ?�B����./��֪F���zj\�D��xm��i8rY�n҃U�,F�_�<3�����h��v#�-ʾ(�y��_C��f��<E����\�d���"�������5�^��_P3틻�Y��^��5�����)�����o���ޯrt�����1��
c�B�b��� 3dE�=		�b9@<��g�~���ރQy$yݻ	�ۿ���L��$��O�M�dP&��%��O1N;~vu5��j�!�No	Y֔Yf=�Է�3���>
���V��b����A<�
�D�
2����K׼/��[���z߀GfH]r�OݕQ�+���j�����N�m�?
޷f����]�==<"v��4c�P»ƭ��ߓ8�a�:�Ǵ��ݓ��OǢlS�ܧXX�^�_]���4\��#�3���Nb���8
�T�KN��;�3�"B����z������㼾=._!�i�����d��io&~���Rw�;1|��})��+��달ѵM�K�kQ��F�'���������z��7�i�y�����(�i-N�Y�_�yT�����|P��|YD��J��!�t�D��>�����wo�B9���3H�ظ����VV�<�>2���Ƴ����kG�T<Z�01	���)tf��N����)�si��c�+�g���e�eVM��B��&)m�N\R�����y�-I���t�h�fWqu�x��,��EN�pǊ(V����;��/�Y���~�6TT#�e
����Rb���-L��Y�VڻwH���Į�CA�+���3ɍ{=;�a�WW1���M��q������ѩ!r�f�˿B;�� 4��Ҥ�m�����I��Տ��zv�`���(��V�Ӓ4CS��1��{�ݗ�Շ]������ ��ƭ�]�'1���0����
i铵�܈|4��Z��%9�tO����~=�pE���T���G�N5��rk�dk������{�b���r��L�|�Nz�ņ�^�B���ʝ��ȋ�A<7�	3q���y�7I��c��Ӵ3� |�)}�N"7�ň�؀ ��ny3�tRW1���~|3�_���i�x��Z+C�Peu��i~�w-�*-8<<|u�y5T�N��7̓NY�Cv�x�g�=ұ�q���bp�V������7���Waۑ��}F��k�A\�x��/�c�Q*�ͣV�Q�/ 'P
����㠐����{m�^
��l|�|�
բ��q��3�8�����[�v��C�gV"�`[Z1XY&[.b��7Q/P�?
L��"�X�'��$>Pu?d� 9���g�Fh7Y�:���ȆA1�����U:���-�ك�L�{�w�S��`	Y�T�y}
�B��&�N"� �Q���W�(��㍺[�=Y3��4��3�Ԅ��JE9�K��#k����;C���:�����<֞���!_�m@(Ca�w�
a�	�_L���O�A{����;1�={1�w�V�H�o�5'.���C�v}fn@���=�8<� n�uA�K��n�O$�z��z+�`{����*�0ۥ݇������]������&���EvMQJ���=?S���:�������S�Q?�׸��|$�p#1��dt#�5��k��r���'r�Z7u���V���^���`���Z��|�,Wv5B��5�&�g3�L�I�s�����]������������EX21'~b,ܚ|��xSe�\�4�z:���R��, ���3#�	�о�9e���d�p�ܿ黈+�(��"�S��-� �Z��%wu�W���7ߟ�t�	���{�vO�V���iNiM)��@��Ȕ��57�*�:�)`ς��|r�21����2�����;��t)2��@}�ʳ�de( ^��f�P� �(��u���ӑx�o��n��qͦ5�\U�{������G���m�� %��Z�T4�R���ni�3�(K�C�+��4�B��܁Lw���@Ђ� eaR�O�KC-�Έv���"�d,�m���]<�w�C����ּ�?f@�[�u�piF��1Ľv���%��
Q.�tg�`N�GA>�o�����������%���/B��R�fnY�a�S�:pm���3~��S�r�nя]D�^>c0�Ȅ����D��KW����+�{O,ɪ�X��@Ѝ� �ԠH	�ͺ��D˟�D\QZ�����#��k�ܰI�̵���̴�@�3%��)���T�:��I��0�<�ym�T@W�/X���Q#ʱ����Z)>B�D�١�1�{]Rr���Y�[�����l�0X�B�x���b�&����8���iQT?�o��3�=b{�a!���X��m�}0��������sE�9����P��[�	~����"'kv':_!\�D�O�� �������zps,��6T���I|!����.����W5�4�|�n����I~ixm�� ���� �;d���eVH��%����"$Q(�����N�!Uσe��M-���Q,d��WM'�u�#���4*5�w>���𠨪 ��_�|
�D��r�K��ȳ��rc*Ŕ���lVk==��)w���Y1wd�7yun�i�8��7�5�f��{3����M�O}�Xy�i<��`ñ�H�\�=~2w��^_\T	���.��y
*��K�D�A���:��;���E���׈k��b��.x���CWw�xyy%���@�عqyY�x����2ň3!����}>-\����\`���o_���Iq����� �a�(׆ѽ	s���=����ܫ��'8��_��w������t�n)f�ƭ����a����h1F*��VM�P�j��;T�X��BY�d���hok�l;��9�1�3}�_�R���6�zyUL�R�܋ �t�>�����7\#M![���Q�6��뗇�W-�/���<@�ë��m����G�|f׾tJ,#�;�=B��Z�;Q����t��f»㥀-��].8�Y�;���"���������]o�/�,Fa��w�b��7\DP�h��X/���m����;�����J:B.�8��*�=���SP��ŞL8{�d���������sD	�j8�pc%��i�ɺ�<�$�x����Qe���&YYyU>s���_f���A��L:^��o��/��gqT2љj�0�X�������l���E�V�vg�y�Y*��P�U��]���q��\����OӜ -�Bk͡���d6r��,I���"˻���/F�C���R%p���5c�7��g�ׂ�H��� 9��g���R��n�-���B����O������4�▣{�c�!�מ���l�@�J��J���&��g��GuuƳA_��6錨�MA��}؜�~A�������t�O�ƙڱ���#��$P^����]ҸN�D:[Z,f=��y��|Z®�ambmm�Y�F;a3��B����n���/
�Iկ��47n�<(�|�OY�et�6s��3M�G=lz�>F �~y)�S
���Ƒ!�aH-�׈9��L�5��9��(��૏��o1��hS�Ce���ȎJ����v"�Ƀ���Z�<�_f6�@�n��-��P���_�h���|[�Ҵ��7�;\��^��_�ǒ͏�O#O�鵿t�ڟ߫簎��^@���sZ��v!�L4�Z~��	m�t��X��8.�ԏ2H������dh3�:�*��tk�/HΧ�FI��X�K��uƺ�W��$b��"�Zg���^1�b�)��-�ҁm���P�	,5!Z��Y4Dp�h3����m��VM�f�K�8�v�Y��c�Ŧ�6O��n[�h{�Hq&
� m���Y�L��$����ŋ>��5;h�W�����i��;m��{�N��Sn�E��ܽ=Q�FZ	Q1���53>\��ghdihȄ+�>�~\�٭x���I�H�zJ%�6OW0�i��,>�X$%/�$'�����?�����Y��T�rЙ�l�,�!~ �[4������!��^Cp뗵)AV!"i�w�#�T>�V��T�N���%v^m��Ž&R���N>?p��5L����q����k$*��� ��,V��p���ϟ&6~(tD�/U�@��$�DC>n��z�2#��gD�n&VI`��ݗ�]��Ǭ�i�-���4�����K���e�p�r!�?ƃ|1�a���{�/=�J�keۼ�~�!�[�q�|5�^�B�@$�8�t�-u���N���k�N�1����u���= Y�+���� �@�*H�._)P�h6@��mb�OHF�FUI���VQ�J�Cz����W|�����ɰ,�	?w�z��(o<* �`~��ۗP���>;��L��V�-+�+��8l=9;����kk�$�i�~��xtZֶ0�OG�,�$\��\��/5Ǘ#�D�R���A���d���˿�-�.����_p�͹u��(�d���R��>���������8���hރ�J11.Le��t�,��p̬a�O�T}����K���0�qƧZ����,�))�nM�=�uA����̏���*ﯰ9�����GCD�\Z-�8��s���Lި�v�Z]]D�Ty����(�O8S5 ��p�HW���G{#�<��ٱ�զW������8}�	Y�t��=��ZDp� rb��Hpön�}T���J�.w�Za�yc�Ϛ���G��ddmb¶7O7�or��U�}@� ����+�*;-G����?� ��_�q��t��b{���%�@��!��MF�߅Ө5t���I�@�H�lh
V������*r�~w�6�t�.����41#x\�G����E_���e�!�J�hD�e�j����Ed�x�Z~y�V��<M���5*��Ⓣ+�;>.��|�^DS
�I"_D(33�u��|��w�H�~Ǵ=�H-�ը�@�� R�Ռ�+�z9;s���b�?r���rso��� fdԙ{@F�o;��$���1꭛�B�!�:������$wZw�
	Y�gt�)OK�[Lp8_.2�d�ǪY��bS�j](b/w��t�s�M��aHC�����8i�w��cu�7s0k�˔zin͓�;��
�=�ӝa����Ҝ��2&��PƇ��hŠ��)�Z)�t�t�c���X�e{7� /Of�rǩu��� (	ܓT�8?���uK�-Jb����J��L��R�_�����} _0H��d�ޞ^��J������ZHo	I�w���A82����'� �-WW>���!�ԟ�>/�.���Ӫ�Y��N"�{P �{��'�~���0��v���}�|��S�q,jw$w����(i͜�,�2ڬ㡀d�T�̓�Θ�*t,	=��3N�,sO�D�k���N,9�Ν+MoHs�ϙ/���~���EC�Yϻ�d��[-܅pà����!���ә��fyḴ�u�o�Aa�W-�mG����Ag�C��\B�z��}#�[��:�Lm7�Y���Ua��Z϶k�:<�;JJ��dK�MOU�+�B4��}�ɟ
<���W�C�^f�B�/2%�;��a�}����B�D��j6����.�(X�3���R��	k{��l�,K��7KezLLL���4o�a�cY��2��A��Dy��hjh�z��Ȭ������*�0{�H�~�N)`�
�����ek�PYsC�&�L*��f�y�X���� h�E�zDߖt�3�?�h���sv�vo���I_���{H�nka��`�D3��`�`f�?ՁI'��	����\��&�B�r��M�����ex����o���G'���=�ث����FS1���� i�^A"��+���vMIc�\�[=��y��'z{�[�˪�|`c
���M]��US��j=j7�N[���pC��׮Օ�k�:�߸m��Uò�t[˿
t��%��ܓ��3(R�Z�_�ǥݢ�|/�xh��q쟚�=cƵ�fϫ��ΫH�x5-���c�(��Jh �Ճ��hG�}y�=��n�m�v��\s����
��Q�$ aM��({M*���W"^*����L?K}QpYv�M�>���x �Ab�7l׬[��'Թ��n�KZ�sA�����Wy� �s���w5k&us��Z"����4��hz��S
#qa�HL�{fYY���ks��0��դ#~@�j= �!YrBޚ��#�G&�-A���?�g� K���E2��S�zvy�zd­�1�w�S��L����z���rlj�c�z�~���,�m���d���h�1����n��3NJ�o@�k����'p�{�:��r������-�X>�gR[Hew�WΧ;Y��k��=D�^�kc�#,�D��ƨ*,�H�p��<P("���Q��q�\Ut�#�{�U���\s���wD�jW1j�E�UF�wv�o{7OE��%Y���*(���I����L3������8��//�b��11�'Q�to�^�?�y�lig8�"��zDd��8I[?\ֺ����b؁f�Y�y�}�Pʃpp�����
�_Q��x^yI#��}	P��%_���	����~��8�^�ɸ���Ǆ��{`��%<���43Y�Uh"O	˷�C̣�bh�R�c���[��գ���'ŉH��I��{��ᨍ�<��Ť8\������Q�s��[��^|j��~Q����/M�����8*�%D�i#Z���%��ě�/m�&K��l� ���:9��������/��@-�<ȍ��I_6 d�h��F�<�1<��#�� ����K��Ǯ��i�4nҀB�|\���,%�O]M��D���j���e���1{%�J�<����F�����K���W�}ͳ�����*]��T$�Z^��*�Y�azb�6 r�� `�W��1e?�&̢�>��2�#f�
�`I�^!S������]����8s{�r��3U�ٗ�����A!$ϓe���_}k����`�q�D�K��o�"�)�	�^���*���5�_��lY�=r�<Ƈ3�)A̗=u�$8�����L�C)\A%	֮O�.��Gd(u׼QS�.��(3���T��F+&)H�.���H��`���=��7�~�<2�c��%"8��U��[���/��2s��:�ߜ:Կ�YoѾu���J�T�����_'	7վ�����G������,��]* ҇���k~���BM��6��͈�6��#w�\�w�tfG6���"�B����V�[�c1�%�p$I�r��n��'��R��7��m9H&-�̋���N!����I���y`�v�1��њy�y���1*�,tu���ο�2T��ݵ�\�/A�׵D|
T�Cق҉.��'��A���J���M���ϭw��������3r�N�8;���Z> l�L=�nrɦ+ϪCA=3!Y�7�����uD�w<:{��i�)��Vd�<�vj����D�~Z�tՋ���ҙ3�b�@��X�8J$ �b^B��V�����G���=Z%l��Jp�1ɨ��ŕ�����,дDN���Y�xG@����c1r#��:=����Z�4�G��}���f$�ro;�]\D@v��'mF��!R��_<�\�Ʉ2W���Yx6��3��Z0�"������73�M�H.�m�3��R�F����W�K��K��7+N"��%|=��5%Ѯ\��������]��0���T͖��R#ڗ��=)���	�͝0�`�5ޭy�C��N���BZ#�N,���̿ު�8�Ǯ�yQ�'_Rs(q��H0��	��Ө�>�o��G�P>j�G��̩���4":�.��C���K��iI��Dّ1�x�)�h(�l�p�@L��`7A46�OI����G�.!"J�����ih;E�v;\qTHUS��:��1�["~�X!AK3��������(N����I	rt�#���vZ@���̡΂��K�j�����*u�z�~ �W�ẔI��O=�4���?==��]w�wG}~������#�'?�c�Ł�o\���J��kn��o�U�&n���$Sr{�v,�v�%7�}Ծ���9�4�Nٴ&�U�]'�P:��i*�zۨ��ѧ-e�C?m����%$__�`x���gMm-䍗F���o1�)\h*������JKD6*U��:-���D�������j��#���`>�C�S{O���E�'z,��/���&����5��:B�L����L<�Q"�&LK|Bg�^�-ؾGp�\�K���B|��6�9�E�G#�.u���^b`����~g��K�L��K�}�ȣ��=UˁzV�j�Z�H����%�aL���Q�����Q{M���~�!!oC�mX�X��w�v�
�'��j=�l���٨9���^N]͟��=<0����IT`X�hP��7: T8�1}���Xj�A��âh8|�C�ZOЯ�AB8��M�Ծ<8�%�����f���gF�$�|ʌC8�lK�4�Z=�S�+����,�׾�)s!���ө�7|����C�")m��Ȥ�k0�U��BT�18�`KT�ޫg������ٱD��{� ���f [4^��?�X$B%.�d}h
t�Rb棕*^�F|H"��bj|����lz��� �0��Hi{CW��%?~s�����B�X��S�v�a(���r�D �70&l�R%cЪ���� ��7@Z\������+H#m��������~�р�:R�z�Fz�u��� '�(>o�$�%2��P#�Y�R�(��so]޸��L (��o�����R���HR
u5i��/?�lGa��-�h�|{4��=���󴲳���@�|}�j=�����A4019��	f`V���S��~_/�I��4%<5���꣠�ގ:�ܹ�JhX:Ʃ��	���&z���2@כ��Wp��" ��^a`���+t#(�f5�����|f<����+�N��)z:}(6�}F�ǡ�\Dg�o�����z&,�\���j,.�lE�X*�&�\2�"bn5P��u�zi��u�L�P�ʘl���L�0R@k��n��C=�ڇ�| ��܉�Ѱt�w�� X��h�n�a^��� �ӏVf���"�>���_5��6��j9��	f���-U�h��_c�6�G�At!�r^�'=�2�4>��7��I"k�w���v[t(���+�JIe�U��G��Ut�.�T�q�/,}��
g�k�w�#�����%��[H�(�2��sc���8�n��+.�+{-	!�,&NƧ��n+}7�AJ��p�+�+�n�ڦ�O7���~N��4U<r�NR�4?�~t�u:������� �M��Q��w����{U��e��,�&�R������pi���]�A��}w���f,�H���uN��~�s��ߤ� ��5�WT��ʜ������1�� Šc���� ���\�������8�U'����KC��#(x�~�E��~ea�����V6�[�N/?җ"�a,�C���Q�~4�����cW$�,��0��}b�f�v���>���s)A1p�[��_�1X� ���s���~�p�J�!;-�����+�y�)ڞ�B���y{~�Ʌ�'k���~�|�tN�J7j�M@�M6Y��NGȱ���5���r��?5Ӟ�m�t�d�my��Ai+��\b#/r;�Fj#�Fx��a
�Ȟ��B(B_��<K*��p�=J��&��&~� ~�l�k�-�^`� �Ҙ�߮�[}�M.��o01�Сh��k����+�z����9M�S�N�7ǘ\]ǩ�1%��7Yu>�N߈G�
�.�����-8 ��������'�f.E�A6O�m%r=�\�l}�Vb�PX5��q!�%�4FR�KA~����z���;��|�g!�--M�ߦ��(
b�G�FM����P@�M��N����۝�=U'�{����Do�R��q�NѢ� �6&�)r"�����1�+���n�4Ͼ����J���8
�a��{
�-�0����#���F��(���\��eī�J9�8m��t�Ukń�?Ց͆:V�-zI1�� ql����+H���$��Ani\8r�@7��5s���<
����ڌ<�����%^[�O?����i㫁�ry�W8�Ȉ�Rc�jv1X	�l�!q��O���
 �������8��H�(��E����}��릈|+�����zFA�fZW�$�!��+0�k �2PO�l���5����Wa?N��6�R�F_��t���:��,B�]3}�ᧈ��c 4g �'�v�|#�9.�������y( -��'vW�M�M�6�G�	'��S١��Оt@�0y���~Fǡ��qo3 �>roS����v��LkE�D+[��h:#��AM��v���a��Y�\�?����XIY�����%����K�y�����^0�ϋ9�~���s��Ia9=��K��� ��1�E�P����1F��6��/�긬Ɋ����>Ըꗙ�,��faK�x���*w��O@xSQ]�!�ğ��K򫋫˂{�
;�>Ol��0Uĳ!��ei���."yZJ�S��.8�I��#7��v�OYZ�������dK�4/薧��5L�CkD�8&L��=�[��Qp�
1���A+��N�	��-a�&X�� >hvǒ�D�!���[<�!�ja�1(ՖY"ԋ�.�.��u2�7#V=*SK�ڟ�.s~ь��	Z�ȹ�:�d�H�&&N67�s�&aZ��1M~�ɪּ��)m;e?!v[�Ě緩^޲\��Ô"�L��\t����
��pnM�hS,����w{������m�4@wި���+��5G`pN�G�NIȻ���//*����@�!�~[A���0�bI(�nӾ<__�'L�#Φs�̱o������n�����f�������do�B����<?��R�����GF���0_j�Yh#w2;�qq'ao�#�{�{.�(��R�-���\`2��G]�F%s�/�s��;�W�M���6g( �FT�u����	��[�T��l�ݿ�.�C�W��v��.����--_ؓ� �=�o�a����2IIIh¦�m��ڵ��9��%Zw�l��S�@#.�ZҎ�E�H�^�����l>RHH�,�|��V���2\`��e*�*�`b"���fpO;�o���:LQC�Kw�_5���L�ވ�*��(c��-J���d�p�b��5�����Pi9����媀~�}G�u�ۺg %>1���DC$����
�y4�X��p�F���t��A�ͣ�j�o���M��ûM&�	�H)��b�H)F��^�LCC�l��j<��NY��+{5��b�ɑ�9����wR^<=~�'�6�߈���&��x�JR��n3!NB�0q�h��Wjn��JBB��������^�c�E"","�y",f����|,,,#,lS&���
p��sv�� O-���O�����������#.#�c�V�K�cH4UuUj����PK   W�dW*'�]L  �
     jsons/user_defined.json��ێ�0�_��X��Il�VP�\t���*Uh�M��%6Is�
!޽β��9���g�쉿���L��
�?F*։���Ry���,L05o��-�����p�Թ6+B'�D0�3�aP��4?�H���Nﲻ)ґ��O���#b�9<�#G�91I��<����%]Rge^�?E,T�:+�^�[��Rgɳ��t�L�͎(�^����a���.����]���k� ��%�gR%�geJH�Ѧ̵�7�W���+����*���)�M��X�B2���$���&���}���7t�v�Ӷ<��q�/�W�/���Z���,X��,��_���.P�3 ��P#l֛m��7�[����U�!�M�uؚOu�v%�g����\ޓy����K�Ə�a��x[����3����T� .@�#)�e:B�����R����y� ��K�w�X)�v�j�اȔs3��ݬ6��^��__��|~}��3��������� tz`�7���<W�r#|nç�aۄ�1��O�CZ�@#D[���� 9�`{JC3�v�M\l{=<h�/�;N��0��yڝ~PK   W�dWi���/  ��            ��    cirkitFile.jsonPK   W�dW)<�4I � /           ��8/  images/3f348383-912a-4adc-88a3-03f2846ee105.pngPK   W�dW�Q��� y� /           ���3 images/7a682d23-8f26-4a7d-8a92-f03913074d3f.pngPK   W�dW*'�]L  �
             ���� jsons/user_defined.jsonPK      <  2�   